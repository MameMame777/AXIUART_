`timescale 1ns / 1ps

// AXIUART_Top System Level Test
// Simple test to verify system-level functionality without complex sequences
class axiuart_system_test extends uart_axi4_base_test;
    
    `uvm_component_utils(axiuart_system_test)
    
    function new(string name = "axiuart_system_test", uvm_component parent = null);
        super.new(name, parent);
    endfunction
    
    virtual function void build_phase(uvm_phase phase);
        super.build_phase(phase);
        `uvm_info("SYSTEM_TEST", "AXIUART_Top System test build phase", UVM_LOW)
    endfunction
    
    virtual task run_phase(uvm_phase phase);
        phase.raise_objection(this, "Starting AXIUART system test");
        
        `uvm_info("SYSTEM_TEST", "=== AXIUART_Top System Test Started ===", UVM_LOW)
        
        // Wait for reset deassertion
        wait (uart_axi4_tb_top.dut.rst == 1'b0);
        repeat (10) @(posedge uart_axi4_tb_top.dut.clk);
        
        `uvm_info("SYSTEM_TEST", "Reset deasserted, system initializing", UVM_LOW)
        
        // Monitor system status
        repeat (50) @(posedge uart_axi4_tb_top.dut.clk);
        
        `uvm_info("SYSTEM_TEST", $sformatf("System Status: Ready=%b, Busy=%b, Error=%b", 
                  uart_axi4_tb_top.dut.system_ready,
                  uart_axi4_tb_top.dut.system_busy, 
                  uart_axi4_tb_top.dut.system_error), UVM_LOW)
        
        // Check internal register block is instantiated
        `uvm_info("SYSTEM_TEST", "Checking internal register block accessibility", UVM_LOW)
        
        // Wait for system to stabilize
        repeat (100) @(posedge uart_axi4_tb_top.dut.clk);
        
        `uvm_info("SYSTEM_TEST", "=== AXIUART_Top System Test Completed Successfully ===", UVM_LOW)
        
        phase.drop_objection(this, "AXIUART system test completed");
    endtask
    
    virtual function void final_phase(uvm_phase phase);
        super.final_phase(phase);
        `uvm_info("SYSTEM_TEST", "*** AXIUART SYSTEM TEST PASSED ***", UVM_LOW)
    endfunction

endclass