`timescale 1ns / 1ps

// Enable simulation-only system status signals
`define DEFINE_SIM

import uvm_pkg::*;
import uart_axi4_test_pkg::*;
`include "uvm_macros.svh"

// Top-level testbench for AXIUART_Top system-level verification
module uart_axi4_tb_top;
    
    // Clock and reset
    logic clk;
    logic rst_n;
    
    // System status signals from DUT (simulation only)
    `ifdef DEFINE_SIM
    logic system_ready;
    logic system_busy;
    logic [7:0] system_error;
    logic bridge_enable_state;
    `endif
    
    // Interface instances
    uart_if uart_if_inst(clk, rst_n);
    bridge_status_if status_if(clk);
    // Note: AXIUART_Top uses internal AXI interface, no external AXI connections

    // Optional internal loopback control (disabled by default)
    localparam bit ENABLE_UART_LOOPBACK = 1'b0;

    // Derived simulation guard to accommodate full register campaigns at 115200 baud
    localparam time SIM_TIMEOUT = 400ms;

    // Ensure the RX line idles high until the driver starts toggling it
    initial begin
        uart_if_inst.uart_rx = 1'b1;
    end
    
    // DUT instance - Using complete AXIUART_Top system
    AXIUART_Top #(
        .CLK_FREQ_HZ(125_000_000),
        .BAUD_RATE(115200),
        .AXI_TIMEOUT(1000),
        .UART_OVERSAMPLE(16),
        .RX_FIFO_DEPTH(64),
        .TX_FIFO_DEPTH(64),
        .MAX_LEN(16),
        .REG_BASE_ADDR(32'h0000_1000)
    ) dut (
        .clk(clk),
        .rst(~rst_n),  // RTL expects active-high reset
        
        // UART interface - external connections
        .uart_rx(uart_if_inst.uart_rx),
        .uart_tx(uart_if_inst.uart_tx),
        .uart_rts_n(uart_if_inst.uart_rts_n),   // Request to Send (active low)
        .uart_cts_n(uart_if_inst.uart_cts_n)    // Clear to Send (active low)
        
        // System status outputs (simulation only)
        `ifdef DEFINE_SIM
        ,
        .system_busy(system_busy),      
        .system_error(system_error),     
        .system_ready(system_ready),
        .bridge_enable_state(bridge_enable_state)
        `endif    
    );

    // Bridge status interface wiring
    assign status_if.rst_n = rst_n;
    `ifdef DEFINE_SIM
    assign status_if.bridge_enable = bridge_enable_state;
    assign status_if.bridge_busy = system_busy;
    assign status_if.bridge_error = system_error;
    assign status_if.system_ready = system_ready;
    `else
    assign status_if.bridge_enable = 1'b0;
    assign status_if.bridge_busy = 1'b0;
    assign status_if.bridge_error = 8'h00;
    assign status_if.system_ready = 1'b0;
    `endif
    
    // *** UART Loopback connection (legacy bring-up mode) ***
    // Disabled for full-system verification so the UVM driver controls uart_rx.
    // Set ENABLE_UART_LOOPBACK=1'b1 if a self-loopback is required for standalone debug.
    generate
        if (ENABLE_UART_LOOPBACK) begin : gen_uart_loopback
            always_comb begin
                uart_if_inst.uart_rx = uart_if_inst.uart_tx;
            end
        end
    endgenerate
    
    // Clock generation (50MHz)
    initial begin
        clk = 1'b0;
        forever #10ns clk = ~clk; // 50MHz clock
    end
    
    // Reset generation
    initial begin
        rst_n = 1'b0;
        repeat (5) @(posedge clk);
        rst_n = 1'b1;
        `uvm_info("TB_TOP", "Reset released", UVM_MEDIUM)
    end
    
    // UVM testbench initialization
    initial begin
        // Import the test package to ensure all classes are registered
        import uart_axi4_test_pkg::*;
        
        // Set virtual interfaces in config database
        uvm_config_db#(virtual uart_if)::set(null, "*", "vif", uart_if_inst);
            uvm_config_db#(virtual uart_if)::set(null, "*", "uart_vif", uart_if_inst); // Legacy support
            uvm_config_db#(virtual bridge_status_if)::set(null, "*", "bridge_status_vif", status_if);
            uvm_config_db#(virtual axi4_lite_if)::set(null, "*", "axi_vif", dut.axi_internal);
        // Note: AXIUART_Top uses internal AXI interface - no external AXI interface to set
        
        // Enable waveform dumping
        $dumpfile("uart_axi4_minimal_test.mxd");
        $dumpvars(0, uart_axi4_tb_top);
        `uvm_info("TB_TOP", "Waveform dumping enabled", UVM_MEDIUM)
        
        // Start UVM test
        run_test();
    end
    
    // Timeout mechanism - extended for comprehensive tests
    initial begin
        #(SIM_TIMEOUT);
        `uvm_error("TB_TOP", $sformatf("Test timeout - simulation exceeded %0t", SIM_TIMEOUT))
        $finish;
    end
    
    // Protocol checker instances for additional verification
    
    // UART protocol checker
    uart_protocol_checker uart_checker (
        .clk(clk),
        .rst_n(rst_n),
        .uart_rx(uart_if_inst.uart_rx),
        .uart_tx(uart_if_inst.uart_tx)
    );
    
    // Note: AXI4-Lite protocol checker not applicable since AXIUART_Top uses internal AXI
    
    // Coverage collection
    `ifdef ENABLE_COVERAGE
        initial begin
            // Enable coverage collection at system level
            // $coverage_control(1);  // Commented out - not supported in all simulators
            `uvm_info("TB_TOP", "Coverage collection enabled", UVM_MEDIUM)
        end
    `endif
    
    // Assertion monitoring (temporarily disabled for compilation)
    `ifdef ENABLE_ASSERTIONS_DISABLED
        // Include assertion bind files for AXIUART_Top
        bind dut uart_axi4_assertions uart_axi4_assert_inst (
            .clk(clk),
            .rst_n(rst_n),
            .uart_rx(uart_rx),
            .uart_tx(uart_tx),
            // AXI interface signals - accessing internal interface
            .axi_awaddr(dut.axi_internal.awaddr),
            .axi_awvalid(dut.axi_internal.awvalid),
            .axi_awready(dut.axi_internal.awready),
            .axi_wdata(dut.axi_internal.wdata),
            .axi_wstrb(dut.axi_internal.wstrb),
            .axi_wvalid(dut.axi_internal.wvalid),
            .axi_wready(dut.axi_internal.wready),
            .axi_bresp(dut.axi_internal.bresp),
            .axi_bvalid(dut.axi_internal.bvalid),
            .axi_bready(dut.axi_internal.bready),
            .axi_araddr(dut.axi_internal.araddr),
            .axi_arvalid(dut.axi_internal.arvalid),
            .axi_arready(dut.axi_internal.arready),
            .axi_rdata(dut.axi_internal.rdata),
            .axi_rresp(dut.axi_internal.rresp),
            .axi_rvalid(dut.axi_internal.rvalid),
            .axi_rready(dut.axi_internal.rready),
            // Bridge internal status - accessing through bridge instance
            .bridge_state(dut.uart_bridge_inst.main_state),
            .frame_complete(dut.uart_bridge_inst.frame_parser.frame_valid),
            .crc_valid(dut.uart_bridge_inst.frame_parser.frame_valid && !dut.uart_bridge_inst.frame_parser.frame_error)
        );
    `endif // ENABLE_ASSERTIONS_DISABLED
    
    // Debug and monitoring for AXIUART_Top
    always @(posedge clk) begin
        if (rst_n) begin
            // Monitor critical signals through bridge instance
            if (dut.uart_bridge_inst.frame_parser.frame_valid) begin
                `uvm_info("TB_TOP", $sformatf("Frame parsed: CMD=0x%02X, ADDR=0x%08X", 
                          dut.uart_bridge_inst.frame_parser.cmd, 
                          dut.uart_bridge_inst.frame_parser.addr), UVM_DEBUG)
            end
            
            // Monitor system status (simulation only)
            `ifdef DEFINE_SIM
            if (dut.system_busy) begin
                `uvm_info("TB_TOP", "System busy", UVM_DEBUG)
            end
            
            if (dut.system_error != 0) begin
                `uvm_info("TB_TOP", $sformatf("System error: 0x%02X", dut.system_error), UVM_HIGH)
            end
            `endif
        end
    end
    
    // Performance monitoring
    real start_time, end_time;
    int transaction_count = 0;
    
    always @(posedge uart_if_inst.uart_rx or posedge uart_if_inst.uart_tx) begin
        if (rst_n) begin
            if ($time > 1000) begin // Skip reset period
                if (transaction_count == 0) start_time = $realtime;
                transaction_count++;
                
                if (transaction_count % 100 == 0) begin
                    end_time = $realtime;
                    `uvm_info("TB_TOP", $sformatf("Processed %0d transactions in %.2f ms", 
                              transaction_count, (end_time - start_time) / 1000000.0), UVM_LOW)
                end
            end
        end
    end
    
    // Save coverage database periodically
    `ifdef ENABLE_COVERAGE
        initial begin
            #2ms;
            `uvm_info("TB_TOP", "Coverage database saved", UVM_MEDIUM)
        end
    `endif
    
endmodule

// UART Protocol Checker
module uart_protocol_checker (
    input logic clk,
    input logic rst_n,
    input logic uart_rx,
    input logic uart_tx
);
    
    // Basic UART frame validation
    // Implementation would include timing checks, frame format validation, etc.
    
endmodule