`timescale 1ns / 1ps

// Import protocol constants from test package
import uart_axi4_test_pkg::*;

// IEEE 1800.2 / UVM Best Practice Compliant UART Driver
// Features:
// - Reset-safe: Uses try_next_item() to avoid deadlock during reset
// - Hang-free: Natural termination support with stop_request
// - Baud-dynamic: Reads baud_rate from config dynamically
// - State-machine based: Proper reset handling
class uart_driver extends uvm_driver #(uart_frame_transaction);
    
    `uvm_component_utils(uart_driver)
    
    // Configuration
    uart_axi4_env_config cfg;
    uvm_tlm_analysis_fifo#(uart_frame_transaction) tx_response_fifo;
    uvm_analysis_port #(uart_frame_transaction) tx_request_ap;
    
    // Virtual interface
    virtual uart_if vif;
    
    // Driver state
    typedef enum {RESET, IDLE, DRIVING, WAIT_RESPONSE} driver_state_t;
    driver_state_t state;
    
    // Runtime parameters (updated from config)
    int current_baud_rate;
    int bit_period_ns;
    int post_frame_idle_cycles;
    
    function new(string name = "uart_driver", uvm_component parent = null);
        super.new(name, parent);
        tx_request_ap = new("tx_request_ap", this);
        state = RESET;
    endfunction
    
    virtual function void build_phase(uvm_phase phase);
        super.build_phase(phase);
        
        // Get configuration
        if (!uvm_config_db#(uart_axi4_env_config)::get(this, "", "cfg", cfg)) begin
            `uvm_fatal("UART_DRIVER", "Failed to get configuration object");
        end
        
        // Get virtual interface
        if (!uvm_config_db#(virtual uart_if)::get(this, "", "vif", vif)) begin
            `uvm_fatal("UART_DRIVER", "Failed to get virtual interface");
        end

        // Optional monitor-provided response FIFO
        if (!uvm_config_db#(uvm_tlm_analysis_fifo#(uart_frame_transaction))::get(this, "", "tx_response_fifo", tx_response_fifo)) begin
            tx_response_fifo = null;
            `uvm_info("UART_DRIVER", "Monitor response FIFO not provided", UVM_LOW);
        end
        
        // Initialize runtime parameters from config
        update_baud_parameters();
    endfunction
    
    // Update baud rate parameters from config (dynamic reconfiguration support)
    virtual function void update_baud_parameters();
        if (cfg == null) return;
        
        current_baud_rate = cfg.baud_rate;
        
        // Calculate bit period in nanoseconds
        // bit_period = (1 / baud_rate) / (1ns)
        // Example: 115200 baud = 8680ns per bit
        bit_period_ns = int'(1_000_000_000.0 / real'(current_baud_rate));
        
        // Get idle cycles from config (default to 20 if not set)
        post_frame_idle_cycles = (cfg.max_idle_cycles > 0) ? cfg.max_idle_cycles : 20;
        
        `uvm_info("UART_DRIVER", $sformatf("Baud parameters updated: rate=%0d, bit_period=%0dns, idle_cycles=%0d",
                  current_baud_rate, bit_period_ns, post_frame_idle_cycles), UVM_MEDIUM);
    endfunction
    
    // UVM Cookbook compliant run_phase
    // Reset is handled by test via uart_reset_seq calling vif.reset_dut()
    // Driver assumes reset already completed when transactions begin
    virtual task run_phase(uvm_phase phase);
        super.run_phase(phase);  // MUST: UVM 1800.2 - Preserve parent objection management and parallel process initialization
        
        begin : run_phase_body
            uart_frame_transaction req;
            
            // Initialize interface signals
            initialize_interface();
            
            `uvm_info("UART_DRIVER", $sformatf("[OK] %s run_phase START (phase=%s)", get_full_name(), phase.get_name()), UVM_LOW);
            `uvm_info("UART_DRIVER", "Run phase started - ready for transactions", UVM_LOW);
            
            // Simple forever loop (UVM Cookbook pattern)
            // No reset handling - test controls reset via sequence
            forever begin
            // Blocking get (IEEE 1800.2 / UVM Cookbook standard)
            `uvm_info("UART_DRIVER", "[DIAGNOSTIC] About to call get_next_item()...", UVM_LOW);
            seq_item_port.get_next_item(req);
            `uvm_info("UART_DRIVER", $sformatf("[OK] Got item of type %s", req.get_type_name()), UVM_LOW);
            
            `uvm_info("UART_DRIVER", $sformatf("Got transaction: CMD=0x%02X ADDR=0x%08X", 
                      req.cmd, req.addr), UVM_MEDIUM);
            
            // Update baud parameters (dynamic support)
            update_baud_parameters();
            
            // State transition
            state = DRIVING;
            
            // Execute transaction
            drive_transaction(req);
            
            // Completion notification (IEEE 1800.2 required)
            `uvm_info("UART_DRIVER", "[CRITICAL_DEBUG] BEFORE item_done() call", UVM_LOW);
            seq_item_port.item_done();
            `uvm_info("UART_DRIVER", "[CRITICAL_DEBUG] AFTER item_done() call", UVM_LOW);
            
            // Post-frame idle (DUT requirement) - skip for reset transactions
            if (!req.is_reset) begin
                apply_post_frame_idle();
            end else begin
                `uvm_info("UART_DRIVER", "Reset transaction - skipping post-frame idle", UVM_HIGH);
            end
            
            `uvm_info("UART_DRIVER", "Transaction completed", UVM_HIGH);
            
            // No objection check needed - driver runs until simulation ends
            // UVM phase mechanism handles proper termination automatically
        end
        
        `uvm_info("UART_DRIVER", "Run phase completed gracefully", UVM_LOW);
        end : run_phase_body
    endtask
    
    // Initialize interface signals
    virtual task initialize_interface();
        vif.uart_rx = 1'b1;    // Idle state (high)
        vif.uart_cts_n = 1'b0; // CTS asserted (ready to receive)
        `uvm_info("UART_DRIVER", "Interface initialized: RX=1 CTS_N=0", UVM_HIGH);
    endtask
    
    // Handle reset transaction (driver-controlled reset via clocking block)
    virtual task handle_reset_transaction(uart_frame_transaction tr);
        `uvm_info("UART_DRIVER", $sformatf("Executing reset transaction: %0d cycles", tr.reset_cycles), UVM_MEDIUM);
        
        // Assert reset (synchronous, active-high)
        vif.driver_cb.rst <= 1'b1;
        vif.driver_cb.rst_n <= 1'b0;
        
        // Hold reset for specified cycles using direct clock edge (not clocking block)
        // This ensures reset works even if clocking block has special reset behavior
        repeat(tr.reset_cycles) @(posedge vif.clk);
        
        // De-assert reset
        @(posedge vif.clk);  // Use direct clock edge - driver_cb may hang if clock stops
        vif.driver_cb.rst <= 1'b0;
        vif.driver_cb.rst_n <= 1'b1;
        
        // Small stabilization delay after reset release
        repeat(5) @(posedge vif.clk);
        
        `uvm_info("UART_DRIVER", "Reset transaction completed", UVM_MEDIUM);
    endtask
    
    // Handle reset event
    virtual task handle_reset();
        if (state != RESET) begin
            `uvm_info("UART_DRIVER", "Reset detected - entering RESET state", UVM_MEDIUM);
            state = RESET;
        end
        
        // Reinitialize interface
        initialize_interface();
        
        // Wait for reset de-assertion (edge-sensitive)
        @(negedge vif.rst);
        
        // Small delay after reset release
        repeat(5) @(posedge vif.clk);
        
        `uvm_info("UART_DRIVER", "Reset de-asserted - returning to IDLE", UVM_MEDIUM);
    endtask
    
    // Drive complete transaction
    virtual task drive_transaction(uart_frame_transaction tr);
        // Check if this is a reset transaction
        if (tr.is_reset) begin
            handle_reset_transaction(tr);
            // No item_done() here - the forever loop handles it after this task returns
            // Early return skips send_frame/collect_response only
            return;
        end
        
        // Check RTS before driving (hardware flow control)
        // RTS is active-low: 1'b0 = ready to receive, 1'b1 = not ready
        `uvm_info("UART_DRIVER", $sformatf("[RTS_CHECK] uart_rts_n=%b before send_frame", vif.uart_rts_n), UVM_LOW);
        
        if (vif.uart_rts_n == 1'b1) begin
            int timeout_cycles = 1000;
            `uvm_warning("UART_DRIVER", $sformatf("RTS de-asserted (uart_rts_n=1) - DUT not ready, waiting (max %0d cycles)...", timeout_cycles));
            
            // Clock-synchronous wait with timeout
            for (int i = 0; i < timeout_cycles; i++) begin
                @(posedge vif.clk);
                if (vif.uart_rts_n == 1'b0) begin
                    `uvm_info("UART_DRIVER", $sformatf("[RTS_RECOVERED] RTS asserted after %0d cycles", i), UVM_LOW);
                    break;
                end
            end
            
            // Final check after timeout
            if (vif.uart_rts_n == 1'b1) begin
                `uvm_error("UART_DRIVER", $sformatf("[RTS_TIMEOUT] RTS still de-asserted after %0d cycles - aborting transaction", timeout_cycles));
                return;  // Abort transaction
            end
        end else begin
            `uvm_info("UART_DRIVER", "[RTS_READY] RTS asserted (uart_rts_n=0) - proceeding with send_frame", UVM_LOW);
        end
        
        // Send frame
        send_frame(tr);
        
        // Handle response if needed
        if (tx_response_fifo != null && !should_skip_response(tr)) begin
            collect_response(tr);
        end
    endtask
    
    // Check if response should be skipped
    virtual function bit should_skip_response(uart_frame_transaction tr);
        // RESET command has no response
        if (tr.cmd == 8'hFF) return 1;
        
        // Baud rate configuration has no response (baud mismatch)
        if (tr.is_write && (tr.addr == 32'h00001008)) return 1;
        
        return 0;
    endfunction
    
    // Send complete UART frame
    virtual task send_frame(uart_frame_transaction tr);
        `uvm_info("UART_DRIVER", $sformatf("Sending frame: SOF=0x%02X CMD=0x%02X ADDR=0x%08X", 
                  SOF_HOST_TO_DEVICE, tr.cmd, tr.addr), UVM_HIGH);
        
        // SOF
        send_uart_byte(SOF_HOST_TO_DEVICE);
        
        // CMD
        send_uart_byte(tr.cmd);
        
        // ADDR (little-endian, 4 bytes)
        send_uart_byte(tr.addr[7:0]);
        send_uart_byte(tr.addr[15:8]);
        send_uart_byte(tr.addr[23:16]);
        send_uart_byte(tr.addr[31:24]);
        
        // DATA (if write command)
        if (tr.cmd[7] == 0 && tr.data.size() > 0) begin
            for (int i = 0; i < tr.data.size(); i++) begin
                send_uart_byte(tr.data[i]);
            end
        end
        
        // CRC (simplified - XOR of CMD and ADDR[7:0])
        send_uart_byte(tr.cmd ^ tr.addr[7:0]);
        
        `uvm_info("UART_DRIVER", "Frame transmission complete", UVM_HIGH);
    endtask
    
    // Send single UART byte (8N1 format) - CLOCK SYNCHRONIZED
    virtual task send_uart_byte(logic [7:0] data);
        int clocks_per_bit;
        
        // Calculate clocks needed per UART bit (convert ns to clock cycles)
        clocks_per_bit = bit_period_ns / 1000; // Assume 1MHz clock (1000ns period)
        if (clocks_per_bit < 1) clocks_per_bit = 1;
        
        // Start bit (low)
        vif.uart_rx = 1'b0;
        repeat (clocks_per_bit) @(posedge vif.clk);
        
        // Data bits (LSB first)
        for (int i = 0; i < 8; i++) begin
            vif.uart_rx = data[i];
            repeat (clocks_per_bit) @(posedge vif.clk);
        end
        
        // Stop bit (high)
        vif.uart_rx = 1'b1;
        repeat (clocks_per_bit) @(posedge vif.clk);
    endtask
    
    // Apply post-frame idle period (critical for DUT idle_cnt)
    virtual task apply_post_frame_idle();
        // Return to idle state
        vif.uart_rx = 1'b1;
        
        // Wait specified idle cycles (allows DUT idle counter to increment)
        repeat(post_frame_idle_cycles) @(posedge vif.clk);
        
        `uvm_info("UART_DRIVER", $sformatf("Post-frame idle applied: %0d cycles", post_frame_idle_cycles), UVM_HIGH);
    endtask
    
    // Collect response from monitor FIFO with timeout
    virtual task collect_response(uart_frame_transaction req);
        uart_frame_transaction rsp;
        bit got_response;
        time timeout_ns;
        
        timeout_ns = cfg.frame_timeout_ns * 4; // Conservative timeout
        got_response = 0;
        
        fork
            begin
                tx_response_fifo.get(rsp);
                got_response = 1;
            end
            begin
                #timeout_ns;
            end
        join_any
        disable fork;
        
        if (got_response) begin
            `uvm_info("UART_DRIVER", $sformatf("Response received: STATUS=0x%02X", rsp.cmd), UVM_MEDIUM);
            req.response_status = rsp.cmd;
            req.response_received = 1;
            req.timeout_error = 0;
        end else begin
            `uvm_warning("UART_DRIVER", "Response timeout - no frame received from DUT");
            req.response_received = 0;
            req.timeout_error = 1;
            req.response_status = STATUS_TIMEOUT;
        end
    endtask
    
    // Reset handler for mid-transaction reset
    virtual task monitor_reset();
        fork
            forever begin
                @(posedge vif.rst);
                `uvm_info("UART_DRIVER", "Asynchronous reset detected", UVM_HIGH);
                // State will be handled in main loop
            end
        join_none
    endtask

endclass
