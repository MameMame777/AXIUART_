`timescale 1ns / 1ps

// UART Monitor for UART-AXI4 Bridge UVM Testbench
class uart_monitor extends uvm_monitor;
    
    `uvm_component_utils(uart_monitor)
    
    // Configuration
    uart_axi4_env_config cfg;
    
    // Virtual interface
    virtual uart_if vif;
    
    // Analysis port for sending collected transactions
    uvm_analysis_port #(uart_frame_transaction) item_collected_port;
    // Alias for environment compatibility
    uvm_analysis_port #(uart_frame_transaction) analysis_port;
    
    // Coverage collection
    uart_axi4_coverage coverage;
    
    // Internal variables
    bit monitor_enabled = 1;
    localparam int MAX_RX_FRAME_BYTES = 80;
    int unsigned rx_publish_count = 0;
    int unsigned tx_publish_count = 0;
    time last_rx_publish_time = 0;
    time last_tx_publish_time = 0;
    
    // ========================================================================
    // State Management (Class-level for reset_sampling_state support)
    // ========================================================================
    // RX path state
    bit rx_waiting_for_sof;
    int rx_byte_count;
    logic [7:0] rx_collected_bytes[];
    int rx_expected_length;
    
    // TX path state
    bit tx_waiting_for_start;
    int tx_byte_count;
    logic [7:0] tx_collected_bytes[];
    int tx_expected_length;
    
    function new(string name = "uart_monitor", uvm_component parent = null);
        super.new(name, parent);
        item_collected_port = new("item_collected_port", this);
        analysis_port = item_collected_port;  // Alias
        rx_publish_count = 0;
        tx_publish_count = 0;
        last_rx_publish_time = 0;
        last_tx_publish_time = 0;
        
        // Initialize state variables
        rx_waiting_for_sof = 1;
        rx_byte_count = 0;
        rx_expected_length = 0;
        tx_waiting_for_start = 1;
        tx_byte_count = 0;
        tx_expected_length = 0;
    endfunction
    
    virtual function void build_phase(uvm_phase phase);
        super.build_phase(phase);
        
        // Get configuration
        if (!uvm_config_db#(uart_axi4_env_config)::get(this, "", "cfg", cfg)) begin
            `uvm_fatal("UART_MONITOR", "Failed to get configuration object")
        end
        
        // Get virtual interface
        if (!uvm_config_db#(virtual uart_if)::get(this, "", "vif", vif)) begin
            `uvm_fatal("UART_MONITOR", "Failed to get virtual interface")
        end
        
        // Get coverage collector
        if (!uvm_config_db#(uart_axi4_coverage)::get(this, "", "coverage", coverage)) begin
            `uvm_info("UART_MONITOR", "Coverage collector not found - coverage disabled", UVM_LOW)
        end
    endfunction
    
    virtual task run_phase(uvm_phase phase);
        `uvm_info("UART_MONITOR", "=== RUN_PHASE STARTED ===", UVM_LOW)
        `uvm_info("UART_MONITOR", "About to fork monitor tasks", UVM_LOW)
        
        // Initialize collection buffers
        rx_collected_bytes = new[100]; // Max frame size
        tx_collected_bytes = new[100]; // Max frame size
        
        fork
            collect_rx_transactions();
            collect_tx_transactions();
            monitor_rts_cts_signals();  // Add flow control monitoring
        join_none
        `uvm_info("UART_MONITOR", "Monitor tasks forked - run_phase returning", UVM_LOW)
        
        // Monitor runs indefinitely until test drops objection
    endtask
    
    // ========================================================================
    // Helper Task: Wait for Signal Edge with Timeout (Unified Pattern)
    // ========================================================================
    virtual task wait_for_edge_with_timeout(
        ref logic signal,
        input logic target_value,
        input time timeout_ns,
        output bit timeout_occurred
    );
        time start_time = $time;
        timeout_occurred = 0;
        
        // Advance at least 1 clock to avoid blocking at time 0
        @(vif.monitor_cb);
        
        while (signal != target_value) begin
            @(vif.monitor_cb);
            if (($time - start_time) >= timeout_ns) begin
                timeout_occurred = 1;
                return;
            end
        end
    endtask
    
    // ========================================================================
    // Helper Function: Create Error Transaction (Unified Pattern)
    // ========================================================================
    virtual function uart_frame_transaction create_error_transaction(
        uart_direction_t dir,
        uart_monitor_parse_error_e error_kind
    );
        uart_frame_transaction tr;
        tr = uart_frame_transaction::type_id::create(
            (dir == UART_RX) ? "uart_rx_error_tr" : "uart_tx_error_tr"
        );
        tr.direction = dir;
        tr.timestamp = $realtime;
        tr.parse_error_kind = error_kind;
        tr.response_received = 0;
        tr.response_status = (error_kind == PARSE_ERROR_TIMEOUT) ? 
                             STATUS_MONITOR_TIMEOUT : STATUS_MONITOR_PARSE_FAIL;
        tr.crc_valid = 0;
        tr.frame_data = new[0];
        tr.frame_length = 0;
        tr.response_data = new[0];
        return tr;
    endfunction
    
    // ========================================================================
    // Monitor RX path (host to device) - REFACTORED
    // ========================================================================
    virtual task collect_rx_transactions();
        uart_frame_transaction tr;
        logic [7:0] temp_byte;
        bit timeout_occurred;
        time rx_delta;
        time rx_wait_timeout_ns;
        
        forever begin
            `uvm_info("UART_MONITOR_DBG", $sformatf("collect_rx_transactions loop tick at time=%0t monitor_enabled=%0d", $time, monitor_enabled), UVM_HIGH)
            if (!monitor_enabled) begin
                @(vif.monitor_cb);
                continue;
            end
            
            if (rx_waiting_for_sof) begin
                // Wait for UART start bit using unified timeout helper
                rx_wait_timeout_ns = (cfg.frame_timeout_ns > 0) ? cfg.frame_timeout_ns : 10_000_000;
                wait_for_edge_with_timeout(vif.uart_rx, 1'b0, rx_wait_timeout_ns, timeout_occurred);
                
                if (timeout_occurred) begin
                    `uvm_info("UART_MONITOR", $sformatf("RX start bit timeout after %0t ns - publishing timeout transaction", rx_wait_timeout_ns), UVM_MEDIUM)
                    tr = create_error_transaction(UART_RX, PARSE_ERROR_TIMEOUT);
                    rx_publish_count++;
                    rx_delta = (last_rx_publish_time != 0) ? ($time - last_rx_publish_time) : 0;
                    `uvm_info("UART_MONITOR", $sformatf("MONITOR_WRITE RX_TIMEOUT @%0t (#%0d delta=%0t)", $time, rx_publish_count, rx_delta), UVM_LOW)
                    last_rx_publish_time = $time;
                    item_collected_port.write(tr);
                    continue;
                end
                
                collect_uart_rx_byte(temp_byte);
                
                // Check if this is a SOF marker
                if (temp_byte == SOF_HOST_TO_DEVICE || temp_byte == SOF_DEVICE_TO_HOST) begin
                    `uvm_info("UART_MONITOR", $sformatf("SOF detected: 0x%02x - Starting frame collection", temp_byte), UVM_MEDIUM)
                    tr = uart_frame_transaction::type_id::create("uart_rx_tr");
                    rx_collected_bytes[0] = temp_byte;
                    rx_byte_count = 1;
                    rx_waiting_for_sof = 0;
                end else begin
                    `uvm_info("UART_MONITOR", $sformatf("Ignoring non-SOF byte: 0x%02x", temp_byte), UVM_HIGH)
                end
            end else begin
                // Collecting frame bytes after SOF
                rx_wait_timeout_ns = (cfg.byte_time_ns > 0) ? (cfg.byte_time_ns * 20) : 2_000_000; // 20 byte times or 2ms
                wait_for_edge_with_timeout(vif.uart_rx, 1'b0, rx_wait_timeout_ns, timeout_occurred);
                
                if (timeout_occurred) begin
                    `uvm_info("UART_MONITOR", $sformatf("Multi-byte timeout after %0d bytes - frame complete", rx_byte_count), UVM_MEDIUM)
                    // Process the collected bytes as complete frame
                    if (rx_byte_count >= 7) begin
                        logic [7:0] frame_bytes_local[];
                        frame_bytes_local = new[rx_byte_count];
                        for (int i = 0; i < rx_byte_count; i++) begin
                            frame_bytes_local[i] = rx_collected_bytes[i];
                        end
                        
                        if (parse_rx_frame(frame_bytes_local, rx_byte_count, tr)) begin
                            tr.direction = UART_RX;
                            tr.timestamp = $realtime;
                            rx_publish_count++;
                            rx_delta = (last_rx_publish_time != 0) ? ($time - last_rx_publish_time) : 0;
                            `uvm_info("UART_MONITOR", $sformatf("MONITOR_WRITE RX @%0t (#%0d delta=%0t): CMD=0x%02X ADDR=0x%08X len=%0d", 
                                      $time, rx_publish_count, rx_delta, tr.cmd, tr.addr, rx_byte_count), UVM_LOW)
                            last_rx_publish_time = $time;
                            item_collected_port.write(tr);
                            if (coverage != null) coverage.sample_uart_transaction(tr);
                        end
                    end
                    rx_waiting_for_sof = 1;
                    rx_byte_count = 0;
                    continue;
                end
                
                collect_uart_rx_byte(temp_byte);
                rx_collected_bytes[rx_byte_count] = temp_byte;
                rx_byte_count++;
                
                `uvm_info("UART_MONITOR", $sformatf("RX byte[%0d]: 0x%02X", rx_byte_count-1, temp_byte), UVM_DEBUG)
                
                // Debug: Show accumulated frame
                if (rx_byte_count <= 10) begin
                    string frame_str = "";
                    for (int i = 0; i < rx_byte_count; i++) begin
                        frame_str = {frame_str, $sformatf("0x%02X ", rx_collected_bytes[i])};
                    end
                    `uvm_info("UART_MONITOR", $sformatf("Frame so far (%0d bytes): %s", rx_byte_count, frame_str), UVM_MEDIUM)
                end
                
                
                // Check if we have enough bytes for a complete frame
                rx_expected_length = calculate_expected_frame_length(rx_collected_bytes, rx_byte_count);

                if (rx_expected_length > 0 && rx_byte_count >= rx_expected_length) begin
                    logic [7:0] frame_bytes_local[];
                    frame_bytes_local = new[rx_expected_length];
                    for (int i = 0; i < rx_expected_length; i++) begin
                        frame_bytes_local[i] = rx_collected_bytes[i];
                    end

                    if (parse_rx_frame(frame_bytes_local, rx_expected_length, tr)) begin
                        tr.direction = UART_RX;
                        tr.timestamp = $realtime;

                        `uvm_info("UART_MONITOR", $sformatf("Successfully parsed RX frame: CMD=0x%02X, ADDR=0x%08X, bytes=%0d", 
                                  tr.cmd, tr.addr, rx_expected_length), UVM_MEDIUM)

                        // Send to analysis port
                        rx_publish_count++;
                        rx_delta = (last_rx_publish_time != 0) ? ($time - last_rx_publish_time) : 0;
                        `uvm_info("UART_MONITOR",
                            $sformatf("MONITOR_WRITE RX @%0t (#%0d delta=%0t): dir=RX CMD=0x%02X ADDR=0x%08X len=%0d status=0x%02X parse_err=%s crc_ok=%0b ts=%0t",
                                $time, rx_publish_count, rx_delta, tr.cmd, tr.addr, rx_expected_length, tr.response_status,
                                tr.parse_error_kind.name(), tr.crc_valid, tr.timestamp),
                            UVM_LOW)
                        last_rx_publish_time = $time;
                        item_collected_port.write(tr);
                        `uvm_info("UART_MONITOR_FIFO",
                            $sformatf("PUSH dir=RX idx=%0d fifo_conn=%s time=%0t",
                                rx_publish_count,
                                (item_collected_port != null) ? "analysis_port" : "NULL",
                                $time),
                            UVM_DEBUG)

                        // Collect coverage
                        if (coverage != null) begin
                            coverage.sample_uart_transaction(tr);
                        end

                        // Reset to wait for next SOF
                        rx_waiting_for_sof = 1;
                        rx_byte_count = 0;
                    end else begin
                        // Parsing failed - reset to search for next frame
                        `uvm_warning("UART_MONITOR", $sformatf("Failed to parse RX frame with expected length %0d - resetting", rx_expected_length))
                        rx_waiting_for_sof = 1;
                        rx_byte_count = 0;
                    end
                end else if (rx_byte_count > MAX_RX_FRAME_BYTES) begin
                    `uvm_warning("UART_MONITOR", $sformatf("Frame length exceeded monitor limit (%0d > %0d) - resetting to wait for SOF", rx_byte_count, MAX_RX_FRAME_BYTES))
                    rx_waiting_for_sof = 1;
                    rx_byte_count = 0;
                end
            end
        end
    endtask
    
    // ========================================================================
    // Monitor TX path (device to host) - REFACTORED
    // ========================================================================
    virtual task collect_tx_transactions();
        uart_frame_transaction tr;
        logic [7:0] temp_byte;
        bit collect_more;
        int bit_time_cycles;
        int inter_byte_timeout_cycles;
        time tx_delta;
        time tx_wait_timeout_ns;
        bit timeout_occurred;
        
        `uvm_info("UART_MONITOR_TX_DEBUG", "=== ENTERING collect_tx_transactions() - Before forever loop ===", UVM_LOW)
        `uvm_info("UART_MONITOR_TX", "=== COLLECT_TX_TRANSACTIONS TASK STARTED ===", UVM_LOW)
        `uvm_info("UART_MONITOR_TX_DEBUG", "Variables initialized - Entering forever loop", UVM_LOW)
        
        forever begin
            `uvm_info("UART_MONITOR_TX_DEBUG", $sformatf("Forever loop iteration start @%0t - monitor_enabled=%0b", $time, monitor_enabled), UVM_MEDIUM)
            
            if (!monitor_enabled) begin
                @(vif.monitor_cb);
                continue;
            end
            
            // Wait for TX start bit using unified timeout helper
            tx_wait_timeout_ns = (cfg.frame_timeout_ns > 0) ? time'(cfg.frame_timeout_ns * 4) : 10_000_000; // 4x frame timeout or 10ms
            `uvm_info("UART_MONITOR_TX_DEBUG", $sformatf("Waiting for TX start with timeout=%0d ns", tx_wait_timeout_ns), UVM_LOW)
            
            // First wait for idle (high)
            wait_for_edge_with_timeout(vif.uart_tx, 1'b1, tx_wait_timeout_ns, timeout_occurred);
            
            if (timeout_occurred) begin
                `uvm_warning("UART_MONITOR_TX_TIMEOUT", $sformatf("TX idle timeout after %0t ns - publishing timeout transaction", tx_wait_timeout_ns))
                tr = create_error_transaction(UART_TX, PARSE_ERROR_TIMEOUT);
                tx_publish_count++;
                tx_delta = (last_tx_publish_time != 0) ? ($time - last_tx_publish_time) : 0;
                `uvm_info("UART_MONITOR", $sformatf("MONITOR_WRITE TX_TIMEOUT @%0t (#%0d delta=%0t)", $time, tx_publish_count, tx_delta), UVM_LOW)
                last_tx_publish_time = $time;
                item_collected_port.write(tr);
                continue;
            end
            
            // Then wait for falling edge (start bit)
            @(negedge vif.uart_tx);
            `uvm_info("UART_MONITOR_TX", $sformatf("Detected TX start edge at %0t", $time), UVM_LOW)
            
            tr = uart_frame_transaction::type_id::create("uart_tx_tr");
            tx_byte_count = 0;
            tx_expected_length = 0;
            collect_more = 1;

            bit_time_cycles = cfg.clk_freq_hz / cfg.baud_rate;
            if (bit_time_cycles < 1) bit_time_cycles = 1;
            inter_byte_timeout_cycles = bit_time_cycles * (cfg.max_idle_cycles + 12);
            
            // Collect frame bytes
            do begin
                collect_uart_tx_byte(temp_byte);
                tx_collected_bytes[tx_byte_count] = temp_byte;
                tx_byte_count++;

                `uvm_info("UART_MONITOR_TX", $sformatf("Collected TX byte[%0d]=0x%02X", tx_byte_count-1, temp_byte), UVM_MEDIUM)

                tx_expected_length = calculate_expected_tx_frame_length(tx_collected_bytes, tx_byte_count);

                if (tx_expected_length > 0 && tx_byte_count >= tx_expected_length) begin
                    collect_more = 0;
                end else begin
                    bit next_byte_pending = 0;

                    fork : tx_frame_collection
                        begin
                            time tx_idle_wait_start = $time;
                            time tx_idle_timeout_ns = (cfg.byte_time_ns > 0) ? (cfg.byte_time_ns * 20) : 2_000_000;
                            while (vif.monitor_cb.uart_tx != 1'b1) begin
                                @(vif.monitor_cb);
                                if (($time - tx_idle_wait_start) >= tx_idle_timeout_ns) break;
                            end
                            if (vif.monitor_cb.uart_tx == 1'b1) begin
                                @(negedge vif.monitor_cb.uart_tx);
                                next_byte_pending = 1;
                            end else begin
                                next_byte_pending = 0;
                            end
                        end
                        begin
                            repeat (inter_byte_timeout_cycles) @(vif.monitor_cb);
                            next_byte_pending = 0;
                        end
                    join_any
                    disable tx_frame_collection;

                    collect_more = next_byte_pending;
                end

            end while (collect_more && tx_byte_count < 100);
            
            // Store raw frame bytes for downstream consumers
            if (tx_byte_count > 0) begin
                tr.frame_data = new[tx_byte_count];
                for (int i = 0; i < tx_byte_count; i++) begin
                    tr.frame_data[i] = tx_collected_bytes[i];
                end
            end
            tr.frame_length = tx_byte_count;

            // Attempt to parse TX frame to populate status/echo/data fields
            tr.direction = UART_TX;
            tr.timestamp = $realtime;
            tr.parse_error_kind = PARSE_ERROR_NONE;
            tr.monitor_recovered = 0;
            if (!parse_tx_frame(tx_collected_bytes, tx_byte_count, tr)) begin
                tr.response_received = 0;
                tr.response_status = STATUS_MONITOR_PARSE_FAIL;
                tr.crc_valid = 0;
                tr.response_data = new[0];
                `uvm_warning("UART_MONITOR", $sformatf("Failed to parse TX frame (%0d bytes) reason=%s", tx_byte_count, tr.parse_error_kind.name()))
            end else begin
                tr.response_received = 1;
            end

            `uvm_info("UART_MONITOR_TX", $sformatf("TX Frame parsed: len=%0d status=0x%02X parse_err=%s", tx_byte_count, tr.response_status, tr.parse_error_kind.name()), UVM_LOW)

            // Send to analysis port
            tx_publish_count++;
            tx_delta = (last_tx_publish_time != 0) ? ($time - last_tx_publish_time) : 0;
            `uvm_info("UART_MONITOR_DBG",
                $sformatf("DBG MONITOR_TX_PUBLISH: @%0t (#%0d delta=%0t) cmd=0x%02X len=%0d status=0x%02X parse_err=%s crc_ok=%0b ts=%0t",
                    $time, tx_publish_count, tx_delta, tr.cmd, tr.frame_length, tr.response_status,
                    tr.parse_error_kind.name(), tr.crc_valid, tr.timestamp),
                UVM_LOW)
            `uvm_info("UART_MONITOR",
                $sformatf("MONITOR_WRITE TX @%0t (#%0d delta=%0t): dir=TX CMD=0x%02X ADDR=0x%08X len=%0d status=0x%02X parse_err=%s crc_ok=%0b ts=%0t",
                    $time, tx_publish_count, tx_delta, tr.cmd, tr.addr, tr.frame_length, tr.response_status,
                    tr.parse_error_kind.name(), tr.crc_valid, tr.timestamp),
                UVM_LOW)
            `uvm_info("UART_MONITOR_TX_PUBLISH",
                $sformatf("TX publish log: time=%0t idx=%0d len=%0d status=0x%02X parse_err=%s subscribers=%0d",
                    $time, tx_publish_count, tr.frame_length, tr.response_status,
                    tr.parse_error_kind.name(), item_collected_port.size()),
                UVM_DEBUG)
            last_tx_publish_time = $time;
            item_collected_port.write(tr);
            `uvm_info("UART_MONITOR_FIFO",
                $sformatf("PUSH dir=TX idx=%0d fifo_conn=%s time=%0t",
                    tx_publish_count,
                    (item_collected_port != null) ? "analysis_port" : "NULL",
                    $time),
                UVM_DEBUG)
            `uvm_info("UART_MONITOR_DBG", $sformatf("analysis_port.write() done for TX #%0d ts=%0t", tx_publish_count, $time), UVM_LOW)
            
            // Collect coverage
            if (coverage != null) begin
                coverage.sample_uart_response(tr);
            end
        end
    endtask
    
    // Collect single byte from RX line - DSIM-SAFE with clocking block
    virtual task collect_uart_rx_byte(output logic [7:0] data);
        // Sample start bit
        repeat (cfg.bit_time_cycles / 2) @(vif.monitor_cb);  // ← CLOCKING BLOCK
        if (vif.monitor_cb.uart_rx != 1'b0) begin
            `uvm_warning("UART_MONITOR", "RX start bit not low")
        end
        
        // Sample data bits (LSB first)
        for (int i = 0; i < 8; i++) begin
            repeat (cfg.bit_time_cycles) @(vif.monitor_cb);  // ← CLOCKING BLOCK
            data[i] = vif.monitor_cb.uart_rx;  // ← Sample via clocking block
        end
        
        // Sample stop bit
        repeat (cfg.bit_time_cycles) @(vif.monitor_cb);  // ← CLOCKING BLOCK
        if (vif.monitor_cb.uart_rx != 1'b1) begin
            `uvm_warning("UART_MONITOR", "RX stop bit not high")
        end
        
        `uvm_info("UART_MONITOR", $sformatf("RX byte: 0x%02X", data), UVM_DEBUG)
    endtask
    
    // Collect single byte from TX line - DSIM-SAFE with clocking block
    virtual task collect_uart_tx_byte(output logic [7:0] data);
        // Sample start bit midpoint
        repeat (cfg.bit_time_cycles / 2) @(vif.monitor_cb);  // ← CLOCKING BLOCK
        `uvm_info("UART_MONITOR_SAMPLE_DEBUG", 
                  $sformatf("Start bit check @ %0t: uart_tx=%0b", $realtime, vif.monitor_cb.uart_tx), UVM_DEBUG)
        if (vif.monitor_cb.uart_tx != 1'b0) begin
            `uvm_info("UART_MONITOR", "TX start bit timing variation detected", UVM_DEBUG)
        end

        // Advance one full bit period to center of data[0]
        repeat (cfg.bit_time_cycles) @(vif.monitor_cb);  // ← CLOCKING BLOCK
        data[0] = vif.monitor_cb.uart_tx;  // ← Sample via clocking block
        `uvm_info("UART_MONITOR_SAMPLE_DEBUG", 
                  $sformatf("data[0]=%0b @ %0t", data[0], $realtime), UVM_DEBUG)
        `uvm_info("UART_MONITOR", $sformatf("Sampled TX data[%0d]=%0b at %0t", 0, data[0], $realtime), UVM_MEDIUM)

        // Sample remaining data bits at full bit intervals
        for (int i = 1; i < 8; i++) begin
            repeat (cfg.bit_time_cycles) @(vif.monitor_cb);  // ← CLOCKING BLOCK
            data[i] = vif.monitor_cb.uart_tx;  // ← Sample via clocking block
            `uvm_info("UART_MONITOR_SAMPLE_DEBUG", 
                      $sformatf("data[%0d]=%0b @ %0t", i, data[i], $realtime), UVM_DEBUG)
            `uvm_info("UART_MONITOR", $sformatf("Sampled TX data[%0d]=%0b at %0t", i, data[i], $realtime), UVM_MEDIUM)
        end

        // Sample stop bit midpoint
        repeat (cfg.bit_time_cycles) @(vif.monitor_cb);  // ← CLOCKING BLOCK
        if (vif.monitor_cb.uart_tx != 1'b1) begin
            `uvm_info("UART_MONITOR", "TX stop bit timing variation detected", UVM_DEBUG)
        end

        `uvm_info("UART_MONITOR_RESULT_DEBUG", 
                  $sformatf("Collected byte=0x%02X (binary: %08b) @ %0t", data, data, $realtime), UVM_DEBUG)
        `uvm_info("UART_MONITOR", $sformatf("TX byte: 0x%02X", data), UVM_DEBUG)
    endtask
    
    // Parse RX frame (host to device)
    virtual function bit parse_rx_frame(logic [7:0] bytes[], int count, uart_frame_transaction tr);
        logic [7:0] calculated_crc;
        string frame_debug = "";
        
        // Debug: Show complete frame being parsed
        for (int i = 0; i < count; i++) begin
            frame_debug = {frame_debug, $sformatf("0x%02X ", bytes[i])};
        end
        `uvm_info("UART_MONITOR", $sformatf("Parsing RX frame (%0d bytes): %s", count, frame_debug), UVM_MEDIUM)
        
        if (count < 7) begin // Minimum: SOF + CMD + ADDR(4) + CRC = 7 bytes
            `uvm_info("UART_MONITOR", $sformatf("RX frame too short: %0d bytes (need at least 7)", count), UVM_MEDIUM)
            return 0;
        end
        
        // Check SOF
        if (bytes[0] != SOF_HOST_TO_DEVICE) begin
            `uvm_info("UART_MONITOR", $sformatf("Invalid SOF: expected=0x%02X, got=0x%02X", 
                      SOF_HOST_TO_DEVICE, bytes[0]), UVM_MEDIUM)
            return 0;
        end
        
        // Extract fields
        tr.cmd = bytes[1];
        tr.addr = {bytes[5], bytes[4], bytes[3], bytes[2]}; // Little-endian
        
        // Extract data for write commands
        if (!tr.cmd[7]) begin // Write command
            int data_bytes = count - 7; // SOF + CMD + ADDR(4) + CRC
            if (data_bytes > 0) begin
                tr.data = new[data_bytes];
                for (int i = 0; i < data_bytes; i++) begin
                    tr.data[i] = bytes[6 + i];
                end
            end
        end
        
        tr.crc = bytes[count - 1];
        
        // Verify CRC (exclude SOF from CRC calculation) 
        calculated_crc = calculate_frame_crc_from_index(bytes, 1, count - 2);
        tr.crc_valid = (tr.crc == calculated_crc);        `uvm_info("UART_MONITOR", $sformatf("CRC validation: received=0x%02X, calculated=0x%02X, valid=%0b", 
                  tr.crc, calculated_crc, tr.crc_valid), UVM_MEDIUM)
        
        if (!tr.crc_valid) begin
            `uvm_warning("UART_MONITOR", $sformatf("CRC mismatch: expected=0x%02X, got=0x%02X", 
                         calculated_crc, tr.crc))
            // For debugging, let's still return success to see if that helps
            // return 0;
        end
        
        `uvm_info("UART_MONITOR", $sformatf("Successfully parsed frame: CMD=0x%02X, ADDR=0x%08X", tr.cmd, tr.addr), UVM_MEDIUM)
        return 1;
    endfunction
    
    // Calculate expected frame length based on command
    virtual function int calculate_expected_frame_length(logic [7:0] bytes[], int current_count);
        logic [7:0] cmd;
        
        if (current_count < 2) 
            calculate_expected_frame_length = 0; // Need at least SOF + CMD
        else begin
            cmd = bytes[1];
            
            if (cmd[7] == 1) begin
                // Read command: SOF + CMD + ADDR[4] + CRC = 7 bytes
                calculate_expected_frame_length = 7;
            end else begin
                int bytes_per_beat;
                int beats;

                case (cmd[5:4])
                    2'b00: bytes_per_beat = 1; // 8-bit
                    2'b01: bytes_per_beat = 2; // 16-bit
                    2'b10: bytes_per_beat = 4; // 32-bit
                    default: bytes_per_beat = 0; // Reserved/invalid sizing
                endcase

                beats = int'(cmd[3:0]) + 1;

                if (bytes_per_beat == 0) begin
                    calculate_expected_frame_length = 0;
                end else begin
                    // SOF + CMD + ADDR(4) + DATA(beats * bytes_per_beat) + CRC
                    calculate_expected_frame_length = 7 + (beats * bytes_per_beat);
                end
            end
        end
    endfunction

    // Calculate expected TX frame length based on status/command
    virtual function int calculate_expected_tx_frame_length(logic [7:0] bytes[], int current_count);
        logic [7:0] status;
        logic [7:0] cmd;
        int bytes_per_beat;
        int beats;

        if (current_count < 2) begin
            return 0; // Need at least SOF + STATUS
        end

        if (bytes[0] != SOF_DEVICE_TO_HOST) begin
            return 0;
        end

        status = bytes[1];

        // Any non-OK status is a short (4-byte) frame: SOF, STATUS, CMD, CRC
        if (status != STATUS_OK) begin
            return 4;
        end

        if (current_count < 3) begin
            return 0; // Need CMD byte to determine format
        end

        cmd = bytes[2];

        // Successful write response (RW=0) is always 4 bytes
        if (cmd[7] == 1'b0) begin
            return 4;
        end

        // Successful read response includes echoed address and payload data
        case (cmd[5:4])
            2'b00: bytes_per_beat = 1;
            2'b01: bytes_per_beat = 2;
            2'b10: bytes_per_beat = 4;
            default: bytes_per_beat = 0;
        endcase

        beats = int'(cmd[3:0]) + 1;

        if (bytes_per_beat == 0) begin
            return 0;
        end

        // SOF + STATUS + CMD + ADDR(4) + DATA + CRC
        return 8 + (beats * bytes_per_beat);
    endfunction
    
    // Parse TX frame (device to host)
    virtual function bit parse_tx_frame(logic [7:0] bytes[], int count, uart_frame_transaction tr);
        logic [7:0] calculated_crc;
        string frame_debug = "";
        
        // Debug: Show complete frame being parsed
        for (int i = 0; i < count; i++) begin
            frame_debug = {frame_debug, $sformatf("0x%02X ", bytes[i])};
        end
        `uvm_info("UART_MONITOR", $sformatf("Parsing TX frame (%0d bytes): %s", count, frame_debug), UVM_MEDIUM)
        
        tr.parse_error_kind = PARSE_ERROR_NONE;

        if (count < 4) begin // Minimum response: SOF + STATUS + CMD + CRC = 4 bytes
            `uvm_info("UART_MONITOR", $sformatf("TX frame too short: %0d bytes (need at least 4)", count), UVM_MEDIUM)
            tr.parse_error_kind = PARSE_ERROR_LENGTH;
            return 0;
        end
        
        // Check SOF
        if (bytes[0] != SOF_DEVICE_TO_HOST) begin
            `uvm_info("UART_MONITOR", $sformatf("Invalid TX SOF: expected=0x%02X, got=0x%02X", 
                     SOF_DEVICE_TO_HOST, bytes[0]), UVM_MEDIUM)
            tr.parse_error_kind = PARSE_ERROR_SOF_MISMATCH;
            return 0;
        end
        
        // Extract status
        tr.response_status = bytes[1];
        tr.response_received = 1;
        
        // Extract echo back fields for verification
        // Error frame: SOF(1) + STATUS(1) + CMD_ECHO(1) + CRC(1) = 4 bytes minimum
        // Success frame: SOF(1) + STATUS(1) + CMD_ECHO(1) + ADDR(4) + DATA + CRC(1) = 8+ bytes
        if (count >= 4) begin
            tr.cmd = bytes[2];  // CMD_ECHO is always at position 2
            if (count >= 7) begin
                tr.addr = {bytes[6], bytes[5], bytes[4], bytes[3]};
            end
        end
        
        // Extract response data (for reads with OK status)
        if (count > 8 && tr.response_status == STATUS_OK) begin
            int data_bytes = count - 8; // SOF + STATUS + CMD + ADDR(4) + CRC
            tr.response_data = new[data_bytes];
            for (int i = 0; i < data_bytes; i++) begin
                tr.response_data[i] = bytes[7 + i];
            end
        end
        
        tr.crc = bytes[count - 1];
        
        // Verify CRC (exclude SOF from CRC calculation)
        calculated_crc = calculate_frame_crc_from_index(bytes, 1, count - 2);
        tr.crc_valid = (tr.crc == calculated_crc);
        
        `uvm_info("UART_MONITOR", $sformatf("TX CRC validation: received=0x%02X, calculated=0x%02X, valid=%0b", 
                  tr.crc, calculated_crc, tr.crc_valid), UVM_MEDIUM)
        
        if (!tr.crc_valid) begin
            `uvm_warning("UART_MONITOR", $sformatf("TX CRC mismatch: expected=0x%02X, got=0x%02X", 
                         calculated_crc, tr.crc))
            tr.parse_error_kind = PARSE_ERROR_CRC;
            // For debugging, let's still return success
            // return 0;
        end
        
        `uvm_info("UART_MONITOR", $sformatf("Successfully parsed TX frame: STATUS=0x%02X, CMD=0x%02X", tr.response_status, tr.cmd), UVM_MEDIUM)
        return 1;
    endfunction
    
    // Calculate CRC8 for frame verification
    virtual function logic [7:0] calculate_frame_crc(logic [7:0] bytes[], int count);
        logic [7:0] crc = 8'h00;
        
        for (int i = 0; i < count; i++) begin
            crc = crc ^ bytes[i];
            for (int j = 0; j < 8; j++) begin
                if (crc[7]) begin
                    crc = (crc << 1) ^ 8'h07; // CRC8 polynomial
                end else begin
                    crc = crc << 1;
                end
            end
        end
        
        return crc;
    endfunction

    // Calculate CRC8 starting from specific index (excludes SOF)
    virtual function logic [7:0] calculate_frame_crc_from_index(logic [7:0] bytes[], int start_idx, int count);
        logic [7:0] crc = 8'h00;
        logic [7:0] crc_temp;
        
        for (int i = start_idx; i < start_idx + count; i++) begin
            // Match RTL implementation: XOR entire byte first, then process 8 bits
            crc_temp = crc ^ bytes[i];
            
            // Process each bit with polynomial 0x07 (matches RTL calc_crc8_byte)
            if (crc_temp[7]) crc_temp = (crc_temp << 1) ^ 8'h07; else crc_temp = crc_temp << 1;
            if (crc_temp[7]) crc_temp = (crc_temp << 1) ^ 8'h07; else crc_temp = crc_temp << 1;
            if (crc_temp[7]) crc_temp = (crc_temp << 1) ^ 8'h07; else crc_temp = crc_temp << 1;
            if (crc_temp[7]) crc_temp = (crc_temp << 1) ^ 8'h07; else crc_temp = crc_temp << 1;
            if (crc_temp[7]) crc_temp = (crc_temp << 1) ^ 8'h07; else crc_temp = crc_temp << 1;
            if (crc_temp[7]) crc_temp = (crc_temp << 1) ^ 8'h07; else crc_temp = crc_temp << 1;
            if (crc_temp[7]) crc_temp = (crc_temp << 1) ^ 8'h07; else crc_temp = crc_temp << 1;
            if (crc_temp[7]) crc_temp = (crc_temp << 1) ^ 8'h07; else crc_temp = crc_temp << 1;
            
            crc = crc_temp;
        end
        
        return crc;
    endfunction
    
    // Control functions
    virtual function void enable_monitor();
        monitor_enabled = 1;
        `uvm_info("UART_MONITOR", "Monitor enabled", UVM_LOW)
    endfunction
    
    virtual function void disable_monitor();
        monitor_enabled = 0;
        `uvm_info("UART_MONITOR", "Monitor disabled", UVM_LOW)
    endfunction

    // Monitor RTS/CTS flow control signals
    virtual task monitor_rts_cts_signals();
        logic prev_rts_n = 1'b1;
        logic prev_cts_n = 1'b1;
        
        forever begin
            @(vif.monitor_cb);  // ← CLOCKING BLOCK
            
            if (!monitor_enabled) continue;
            
            // Monitor RTS signal changes
            if (vif.uart_rts_n !== prev_rts_n) begin
                `uvm_info("UART_MONITOR", $sformatf("RTS signal changed: %s", 
                          vif.uart_rts_n ? "deasserted (high)" : "asserted (low)"), UVM_MEDIUM);
                prev_rts_n = vif.uart_rts_n;
            end
            
            // Monitor CTS signal changes
            if (vif.uart_cts_n !== prev_cts_n) begin
                `uvm_info("UART_MONITOR", $sformatf("CTS signal changed: %s", 
                          vif.uart_cts_n ? "deasserted (high)" : "asserted (low)"), UVM_MEDIUM);
                prev_cts_n = vif.uart_cts_n;
            end
        end
    endtask

    // Check for flow control violations
    virtual function bit check_flow_control_violation();
        // Check if transmission occurred while CTS was deasserted
        if (vif.uart_cts_n == 1'b1 && vif.uart_tx == 1'b0) begin
            `uvm_error("UART_MONITOR", "Flow control violation: TX transmission while CTS deasserted");
            return 1;
        end
        return 0;
    endfunction

    // ========================================================================
    // Baud rate 切替時の状態リセット (Refactored)
    // ========================================================================
    // CONFIG write 後のゴミデータ（baud rate 不一致期間のサンプリング結果）を破棄
    // Test 側から明示的に呼び出される
    virtual function void reset_sampling_state();
        `uvm_info(get_type_name(), 
            $sformatf("Resetting sampling state @ t=%0t for baud rate change", $time),
            UVM_HIGH)
        
        `uvm_info(get_type_name(), 
            $sformatf("Discarding stale sampling state (published: RX=%0d TX=%0d, buffered: RX=%0d TX=%0d bytes)", 
                      rx_publish_count, tx_publish_count, rx_byte_count, tx_byte_count),
            UVM_MEDIUM)
        
        // Reset RX path state (now class-level variables)
        rx_waiting_for_sof = 1;
        rx_byte_count = 0;
        rx_expected_length = 0;
        if (rx_collected_bytes != null) rx_collected_bytes = new[0];
        
        // Reset TX path state (now class-level variables)
        tx_waiting_for_start = 1;
        tx_byte_count = 0;
        tx_expected_length = 0;
        if (tx_collected_bytes != null) tx_collected_bytes = new[0];
        
        `uvm_info(get_type_name(), 
            "Sampling state reset complete - ready for new baud rate frames",
            UVM_HIGH)
    endfunction

endclass