`timescale 1ns / 1ps

//==============================================================================
// Register Block Comprehensive Test Sequence
// 
// Purpose: Detailed verification of all Register_Block.sv functions
//          that are NOT covered by current high-level UVM tests
//
// Test Categories:
// 1. Individual Register Access Tests
// 2. Address Validation Function Tests  
// 3. Error Condition Tests
// 4. AXI4-Lite Protocol Compliance Tests
// 5. Data Accuracy Verification Tests
//
// Author: UVM Verification Team
// Date: 2025-10-09
// Version: 1.0
//==============================================================================

// This sequence must be included in uart_axi4_test_pkg.sv
class register_block_comprehensive_sequence extends uvm_sequence#(uart_frame_transaction);
    `uvm_object_utils(register_block_comprehensive_sequence)
    
    // Complete register test specification
    typedef struct {
        string name;
        bit [31:0] address;
        bit [31:0] test_data;
        bit [31:0] expected_readback;
        bit expect_error;
        bit is_read_only;
        string description;
    } register_test_t;
    
    register_test_t register_tests[$];
    
    function new(string name = "register_block_comprehensive_sequence");
        super.new(name);
        create_register_tests();
    endfunction
    
    function void create_register_tests();
        register_test_t test;
        
        // === SYSTEM REGISTERS TEST ===
        
        // Test 1: REG_CONTROL (0x1000) - Read/Write 
        test.name = "control_register_test";
        test.address = 32'h0000_1000;
        test.test_data = 32'h12345679; // Test value for control register
        test.expected_readback = 32'h12345679;
        test.expect_error = 0;
        test.is_read_only = 0;
        test.description = "Control register read/write functionality";
        register_tests.push_back(test);
        
        // Test 2: REG_STATUS (0x1004) - Read Only (composite)
        test.name = "status_register_test";
        test.address = 32'h0000_1004;
        test.test_data = 32'hDEADBEEF; // Should be ignored
        test.expected_readback = 32'h0; // Status bits from bridge inputs
        test.expect_error = 0;
        test.is_read_only = 1;
        test.description = "Status register read-only verification";
        register_tests.push_back(test);
        
        // Test 3: REG_CONFIG (0x1008) - Read/Write
        test.name = "config_register_test";
        test.address = 32'h0000_1008;
        test.test_data = 32'hAABBCCDD;
        test.expected_readback = 32'hAABBCCDD;
        test.expect_error = 0;
        test.is_read_only = 0;
        test.description = "Configuration register functionality";
        register_tests.push_back(test);
        
        // Test 4: REG_VERSION (0x101C) - Read Only  
        test.name = "version_register_test";
        test.address = 32'h0000_101C;
        test.test_data = 32'h11111111; // Should be ignored
        test.expected_readback = 32'h00010001; // Fixed version
        test.expect_error = 0;
        test.is_read_only = 1;
        test.description = "Version register read-only verification";
        register_tests.push_back(test);
        
        // === TEST REGISTERS SET ===
        
        // Test 5: REG_TEST_0 (0x1020) - Basic Read/Write
        test.name = "test_register_0";
        test.address = 32'h0000_1020;
        test.test_data = 32'h55AA55AA;
        test.expected_readback = 32'h55AA55AA;
        test.expect_error = 0;
        test.is_read_only = 0;
        test.description = "Test register 0 - basic read/write";
        register_tests.push_back(test);
        
        // Test 6: REG_TEST_1 (0x1024) - Pattern Test
        test.name = "test_register_1";
        test.address = 32'h0000_1024;
        test.test_data = 32'hF0F0F0F0;
        test.expected_readback = 32'hF0F0F0F0;
        test.expect_error = 0;
        test.is_read_only = 0;
        test.description = "Test register 1 - pattern verification";
        register_tests.push_back(test);
        
        // Test 7: REG_TEST_4 (0x1040) - Gap Address Test
        test.name = "test_register_4_gap";
        test.address = 32'h0000_1040;
        test.test_data = 32'h12345678;
        test.expected_readback = 32'h12345678;
        test.expect_error = 0;
        test.is_read_only = 0;
        test.description = "Test register 4 - gap address handling";
        register_tests.push_back(test);
        
        // Test 8: REG_TEST_7 (0x1100) - Extended Range
        test.name = "test_register_7_extended";
        test.address = 32'h0000_1100;
        test.test_data = 32'hFFFFFFFF;
        test.expected_readback = 32'hFFFFFFFF;
        test.expect_error = 0;
        test.is_read_only = 0;
        test.description = "Test register 7 - extended address range";
        register_tests.push_back(test);
        
        // === ERROR CONDITION TESTS ===
        
        // Test 9: Invalid Address (Below Range)
        test.name = "invalid_address_below";
        test.address = 32'h0000_0FFF; // Below BASE_ADDR
        test.test_data = 32'h00000000;
        test.expected_readback = 32'h00000000;
        test.expect_error = 1;
        test.is_read_only = 0;
        test.description = "Invalid address below range - should return error";
        register_tests.push_back(test);
        
        // Test 10: Invalid Address (Above Range)
        test.name = "invalid_address_above";
        test.address = 32'h0000_1200; // Above valid range
        test.test_data = 32'h00000000;
        test.expected_readback = 32'h00000000;
        test.expect_error = 1;
        test.is_read_only = 0;
        test.description = "Invalid address above range - should return error";
        register_tests.push_back(test);
        
        // Test 11: Unaligned Address
        test.name = "unaligned_address";
        test.address = 32'h0000_1001; // Unaligned (should be multiple of 4)
        test.test_data = 32'h00000000;
        test.expected_readback = 32'h00000000;
        test.expect_error = 1;
        test.is_read_only = 0;
        test.description = "Unaligned address - should return error";
        register_tests.push_back(test);
        
        // === BOUNDARY CONDITION TESTS ===
        
        // Test 12: Address at BASE_ADDR boundary
        test.name = "boundary_base_addr";
        test.address = 32'h0000_1000; // Exactly at BASE_ADDR
        test.test_data = 32'hBEEFCAFE;
        test.expected_readback = 32'hBEEFCAFE;
        test.expect_error = 0;
        test.is_read_only = 0;
        test.description = "Boundary test - exact BASE_ADDR";
        register_tests.push_back(test);
        
        `uvm_info("REG_SEQ", $sformatf("Created %0d comprehensive register tests", 
                 register_tests.size()), UVM_MEDIUM)
    endfunction
    
    virtual task body();
        uart_frame_transaction req;
        int test_num = 0;
        int pass_count = 0;
        int fail_count = 0;
        
        `uvm_info("REG_SEQ", "=== Starting Register Block Comprehensive Testing ===", UVM_LOW)
        `uvm_info("REG_SEQ", "Testing ALL register functions missing from current UVM", UVM_LOW)
        
        foreach (register_tests[i]) begin
            test_num++;
            
            `uvm_info("REG_SEQ", $sformatf("Test %0d/%0d: %s", 
                     test_num, register_tests.size(), register_tests[i].name), UVM_MEDIUM)
            `uvm_info("REG_SEQ", $sformatf("Address: 0x%08X, Data: 0x%08X", 
                     register_tests[i].address, register_tests[i].test_data), UVM_MEDIUM)
            `uvm_info("REG_SEQ", $sformatf("Description: %s", register_tests[i].description), UVM_MEDIUM)
            
            // Execute write operation (if not read-only)
            if (!register_tests[i].is_read_only) begin
                execute_register_write(register_tests[i]);
                `uvm_info("REG_SEQ", "✅ Write operation completed", UVM_MEDIUM)
            end
            
            // Execute read operation and verify
            execute_register_read_verify(register_tests[i]);
            `uvm_info("REG_SEQ", "✅ Read operation completed", UVM_MEDIUM)
            pass_count++;
            
            // Delay between tests
            #(5us);
        end
        
        `uvm_info("REG_SEQ", $sformatf("=== Register Testing Complete: %0d PASS, %0d FAIL ===", 
                 pass_count, fail_count), UVM_LOW)
    endtask
    
    // Helper task: Execute register write operation
    virtual task execute_register_write(register_test_t test);
        uart_frame_transaction req;
        
        `uvm_info("REG_SEQ", $sformatf("Writing 0x%08X to address 0x%08X", 
                 test.test_data, test.address), UVM_HIGH)
        
        // Create and send transaction
        req = uart_frame_transaction::type_id::create("write_req");
        start_item(req);
        
        // Set transaction fields directly (not frame_data array)
        req.cmd = 8'h20;  // 32-bit write command
        req.addr = test.address;
        req.data = new[4];
        req.data[0] = test.test_data[7:0];
        req.data[1] = test.test_data[15:8];
        req.data[2] = test.test_data[23:16];
        req.data[3] = test.test_data[31:24];
        
        req.expect_error = test.expect_error;
        finish_item(req);
    endtask
    
    // Helper task: Execute register read and verify
    virtual task execute_register_read_verify(register_test_t test);
        uart_frame_transaction req;
        
        `uvm_info("REG_SEQ", $sformatf("Reading from address 0x%08X, expecting 0x%08X", 
                 test.address, test.expected_readback), UVM_HIGH)
        
        // Create and send transaction
        req = uart_frame_transaction::type_id::create("read_req");
        start_item(req);
        
        // Set transaction fields directly (not frame_data array)
        req.cmd = 8'hA0;  // 32-bit read command
        req.addr = test.address;
        req.data = new[0]; // No data for read operation
        
        req.expect_error = test.expect_error;
        // Note: expected_read_data is handled by the monitor
        finish_item(req);
    endtask
    
endclass : register_block_comprehensive_sequence