`timescale 1ns / 1ps

// Enhanced UART AXI4 Base Test with Mandatory Reporting Standards
// Created: October 10, 2025
// Purpose: Default enhanced reporting for all future UVM tests

class enhanced_uart_axi4_base_test extends uart_axi4_base_test;
    
    `uvm_component_utils(enhanced_uart_axi4_base_test)
    
    function new(string name = "enhanced_uart_axi4_base_test", uvm_component parent = null);
        super.new(name, parent);
    endfunction
    
    // Enhanced build phase with mandatory reporting configuration
    virtual function void build_phase(uvm_phase phase);
        super.build_phase(phase);
        
        // Configure enhanced reporting as default standard
        configure_default_reporting();
        
        `uvm_info("ENHANCED_BASE", "Enhanced UVM reporting configured for all tests", UVM_LOW)
    endfunction
    
    // Mandatory reporting configuration for all tests
    virtual function void configure_default_reporting();
        uvm_report_server server = uvm_report_server::get_server();
        
        // Standard verbosity hierarchy (October 10, 2025 specification)
        this.set_report_verbosity_level_hier(UVM_MEDIUM);
        this.set_report_verbosity_level_hier(UVM_HIGH);
        this.set_report_verbosity_level_hier(UVM_MEDIUM);
        this.set_report_verbosity_level_hier(UVM_LOW);
        this.set_report_verbosity_level_hier(UVM_LOW);
        this.set_report_verbosity_level_hier(UVM_MEDIUM);
        
        // Configure report actions for enhanced analysis
        this.set_report_id_action_hier("*", UVM_DISPLAY | UVM_LOG | UVM_COUNT);
        this.set_report_id_action_hier("ERROR_*", UVM_DISPLAY | UVM_LOG | UVM_COUNT | UVM_EXIT);
        this.set_report_id_action_hier("FATAL_*", UVM_DISPLAY | UVM_LOG | UVM_COUNT | UVM_EXIT);
        
        // Test-specific verbosity optimization
        configure_component_verbosity();
        
        `uvm_info("ENHANCED_REPORTING", "Default enhanced reporting configuration complete", UVM_LOW)
    endfunction
    
    // Component-specific verbosity optimization
    virtual function void configure_component_verbosity();
        // Reduce noise from high-volume components
        this.set_report_verbosity_level_hier(UVM_LOW);
        
        // Enhance critical path visibility
        this.set_report_verbosity_level_hier(UVM_MEDIUM);
        this.set_report_verbosity_level_hier(UVM_MEDIUM);
        
        // Coverage and analysis components
        this.set_report_verbosity_level_hier(UVM_MEDIUM);
        this.set_report_verbosity_level_hier(UVM_HIGH);
        
        `uvm_info("COMPONENT_CONFIG", "Component-specific verbosity configured", UVM_LOW)
    endfunction
    
    // Enhanced connect phase with reporting validation
    virtual function void connect_phase(uvm_phase phase);
        super.connect_phase(phase);
        
        // Validate reporting configuration
        validate_reporting_setup();
    endfunction
    
    // Reporting configuration validation
    virtual function void validate_reporting_setup();
        uvm_report_server server = uvm_report_server::get_server();
        
        `uvm_info("REPORTING_VALIDATION", "Enhanced reporting setup validated", UVM_LOW)
        `uvm_info("REPORTING_CONFIG", $sformatf("Report server: %s", server.get_name()), UVM_MEDIUM)
    endfunction
    
    // Enhanced test startup with reporting announcement
    virtual task run_phase(uvm_phase phase);
        `uvm_info("ENHANCED_TEST_START", 
                 $sformatf("Starting enhanced test: %s with mandatory reporting", get_name()), UVM_LOW)
        
        // Call parent run_phase
        super.run_phase(phase);
        
        `uvm_info("ENHANCED_TEST_COMPLETE", "Enhanced test execution completed", UVM_LOW)
    endtask
    
    // Enhanced final phase with report summary
    virtual function void final_phase(uvm_phase phase);
        super.final_phase(phase);
        
        // Generate enhanced test summary
        generate_enhanced_summary();
    endfunction
    
    // Enhanced test summary generation
    virtual function void generate_enhanced_summary();
        uvm_report_server server = uvm_report_server::get_server();
        
        `uvm_info("ENHANCED_SUMMARY", "=== ENHANCED TEST SUMMARY ===", UVM_LOW)
        `uvm_info("ENHANCED_SUMMARY", $sformatf("Test: %s", get_name()), UVM_LOW)
        `uvm_info("ENHANCED_SUMMARY", "Enhanced reporting features enabled", UVM_LOW)
        `uvm_info("ENHANCED_SUMMARY", "Report analysis ready for PowerShell processing", UVM_LOW)
    endfunction
    
endclass : enhanced_uart_axi4_base_test