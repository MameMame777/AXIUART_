`timescale 1ns / 1ps

// UVM Test Package for UART-AXI4 Bridge
// Contains all UVM components, sequences, tests, and utilities
package uart_axi4_test_pkg;
    
    import uvm_pkg::*;
    `include "uvm_macros.svh"
    
    // UVM Analysis Port Declarations (must be before class definitions)
    `uvm_analysis_imp_decl(_uart)
    `uvm_analysis_imp_decl(_axi)
    `uvm_analysis_imp_decl(_dut)

    // Protocol constants (FIXED BAUD RATE: 115200 bps)
    parameter int CLK_FREQ_HZ = 125_000_000;
    parameter int UART_OVERSAMPLE = 16;
    parameter int BAUD_RATE = 115200;  // FIXED: 115200 bps
    parameter int BIT_TIME_NS = 1_000_000_000 / BAUD_RATE;  // 8680 ns per bit
    parameter int BYTE_TIME_NS = BIT_TIME_NS * 10; // 8 data + 1 start + 1 stop

    // Configuration class (must appear before any component that consumes it)
    `include "../env/uart_axi4_env_config.sv"

    // Transaction direction constants
    typedef enum { UART_RX, UART_TX } uart_direction_t;
    typedef enum { AXI_WRITE, AXI_READ } axi_trans_type_t;
    typedef enum logic [1:0] { AXI_OKAY = 2'b00, AXI_EXOKAY = 2'b01, AXI_SLVERR = 2'b10, AXI_DECERR = 2'b11 } axi_response_t;

    // DUT Transaction Types  
    typedef enum {
        UART_RX_DATA, 
        FRAME_START_DETECTED, 
        FRAME_COMPLETE,
        AXI_WRITE_ADDR,
        AXI_WRITE_DATA, 
        AXI_WRITE_RESP,
        AXI_READ_ADDR,
        AXI_READ_DATA,
        INTERNAL_STATE_CHANGE,
        FIFO_STATUS_CHANGE
    } dut_transaction_type_t;
    
    // Frame constants from protocol specification
    parameter logic [7:0] SOF_HOST_TO_DEVICE = 8'hA5;  // Host to device SOF (corrected to match RTL)
    parameter logic [7:0] SOF_DEVICE_TO_HOST = 8'h5A;  // Device to host SOF (matches RTL Frame_Builder)
    
    // Command constants
    parameter logic [7:0] READ_CMD  = 8'h80;  // Read command (bit 7 = 1)
    parameter logic [7:0] WRITE_CMD = 8'h00;  // Write command (bit 7 = 0)
    
    // Register addresses for testing
    parameter logic [31:0] TEST_REG_ADDR        = 32'h0000_1020;
    parameter logic [31:0] STATUS_REG_ADDR      = 32'h0000_1004;
    parameter logic [31:0] FIFO_STATUS_REG_ADDR = 32'h0000_1018;
    
    // Status codes
    parameter logic [7:0] STATUS_OK         = 8'h00;
    parameter logic [7:0] STATUS_CRC_ERR    = 8'h01;
    parameter logic [7:0] STATUS_CMD_INV    = 8'h02;
    parameter logic [7:0] STATUS_ADDR_ALIGN = 8'h03;
    parameter logic [7:0] STATUS_TIMEOUT    = 8'h04;
    parameter logic [7:0] STATUS_AXI_SLVERR = 8'h05;
    parameter logic [7:0] STATUS_BUSY       = 8'h06;
    parameter logic [7:0] STATUS_LEN_RANGE  = 8'h07;
    parameter logic [7:0] STATUS_MONITOR_PARSE_FAIL = 8'hF0;
    parameter logic [7:0] STATUS_MONITOR_TIMEOUT    = 8'hF1;

    typedef enum logic [2:0] {
        PARSE_ERROR_NONE,
        PARSE_ERROR_SOF_MISMATCH,
        PARSE_ERROR_LENGTH,
        PARSE_ERROR_STOP_BIT,
        PARSE_ERROR_CRC,
        PARSE_ERROR_PAYLOAD,
        PARSE_ERROR_TIMEOUT
    } uart_monitor_parse_error_e;
    
    // Additional enum types for QA-2.1 Enhanced Scoreboard and DUT Monitor  
    // Note: Using existing axi_trans_type_t for transaction types (AXI_READ, AXI_WRITE)
    // Note: Using existing axi_response_t for response types (AXI_OKAY, AXI_EXOKAY, etc.)
    
    // Additional DUT Transaction Types (complementing dut_transaction_type_t)
    typedef enum {
        UART_TX_START,
        UART_TX_COMPLETE,
        FRAME_PARSING_ERROR,
        CRC_CHECK_RESULT
    } additional_dut_transaction_type_t;
    
    // CRC8 calculation function (polynomial 0x07)
    function automatic logic [7:0] calculate_crc8(input logic [7:0] data[], input int length);
        logic [7:0] crc = 8'h00;
        logic [7:0] temp;
        
        for (int i = 0; i < length; i++) begin
            temp = crc ^ data[i];
            for (int j = 0; j < 8; j++) begin
                if (temp[7]) begin
                    temp = (temp << 1) ^ 8'h07;
                end else begin
                    temp = temp << 1;
                end
            end
            crc = temp;
        end
        return crc;
    endfunction
    
    // UART frame transaction class
    class uart_frame_transaction extends uvm_sequence_item;
        
        // Frame fields - standardized naming
        rand logic [7:0]  sof;      // Start of Frame byte
        rand logic [7:0]  cmd;
        logic [31:0] addr;          // CRITICAL: Remove rand to prevent randomization override
        rand logic [7:0]  len;      // Length byte
        logic [7:0]  data[];        // CRITICAL: Remove rand to prevent randomization override
        logic [7:0]       crc;
        
        // Standardized frame fields for compatibility
        rand logic [7:0]  frame_data[];  // Complete frame data including SOF, CMD, ADDR, DATA, CRC
        rand int          frame_length;  // Total frame length in bytes
        
        // Additional frame analysis fields
        logic [7:0] start_delimiter;   // Same as sof but for scoreboard compatibility
        logic [7:0] crc_received;      // CRC received in frame
        logic [7:0] crc_calculated;    // CRC calculated from data
        int data_length;               // Data payload length  
        logic [7:0] payload_data[];    // Payload data array
        
        // Transaction type
        rand bit is_write;
        rand bit auto_increment;
        rand logic [1:0] size;  // 00=8bit, 01=16bit, 10=32bit, 11=reserved
        rand logic [3:0] length; // 0-15 (actual length is length+1)
        
        // Reset transaction fields
        bit is_reset = 0;           // Flag indicating this is a reset transaction
        int reset_cycles = 100;     // Number of clock cycles to hold reset
        
        // Transaction direction and timing
        uart_direction_t direction;
        realtime timestamp;
        bit crc_valid;
        
        // Error injection fields - standardized
        bit force_crc_error = 0;
        bit force_timeout = 0;
        bit corrupt_frame_format = 0;
        bit truncate_frame = 0;
        bit wrong_sof = 0;
        bit error_inject = 0;        // General error injection flag
    bit expect_error = 0;         // Expect an error response from DUT
        bit data_randomization = 0;  // Data randomization control
        
        // Response fields
        logic [7:0] response_status;
        logic [7:0] response_data[];
        bit response_received;
        
        // Coverage support fields (for axiuart_cov_pkg)
        logic [31:0] target_addr;    // Alias for addr
        bit [6:0]    rx_fifo_level;  // FIFO monitoring
        bit [6:0]    tx_fifo_level;  // FIFO monitoring
        bit          parity_error;   // Error flags
        bit          framing_error;
        bit          timeout_error;
        bit [2:0]    parser_state;   // FSM states
        bit [2:0]    axi_state;
    bit [2:0]    frame_type;     // Derived field
    bit [7:0]    crc_result;     // CRC calculation result
    uart_monitor_parse_error_e parse_error_kind;
    bit          monitor_recovered;
        
        // Constraints
        constraint c_valid_size { size inside {2'b00, 2'b01, 2'b10}; }
        constraint c_valid_length { length <= 15; } // Max 16 beats
        // Note: data size constraint removed as data is now non-rand and managed explicitly
        
        `uvm_object_utils_begin(uart_frame_transaction)
            `uvm_field_int(sof, UVM_ALL_ON)
            `uvm_field_int(cmd, UVM_ALL_ON)
            `uvm_field_int(addr, UVM_ALL_ON)
            `uvm_field_int(len, UVM_ALL_ON)
            `uvm_field_array_int(data, UVM_ALL_ON)
            `uvm_field_int(crc, UVM_ALL_ON)
            `uvm_field_array_int(frame_data, UVM_ALL_ON)
            `uvm_field_int(frame_length, UVM_ALL_ON)
            `uvm_field_int(is_write, UVM_ALL_ON)
            `uvm_field_int(auto_increment, UVM_ALL_ON)
            `uvm_field_int(size, UVM_ALL_ON)
            `uvm_field_int(length, UVM_ALL_ON)
            `uvm_field_int(is_reset, UVM_ALL_ON)
            `uvm_field_int(reset_cycles, UVM_ALL_ON)
            `uvm_field_enum(uart_direction_t, direction, UVM_ALL_ON)
            `uvm_field_real(timestamp, UVM_ALL_ON)
            `uvm_field_int(crc_valid, UVM_ALL_ON)
            `uvm_field_int(error_inject, UVM_ALL_ON)
            `uvm_field_int(data_randomization, UVM_ALL_ON)
            `uvm_field_int(expect_error, UVM_ALL_ON)
            `uvm_field_int(response_status, UVM_ALL_ON)
            `uvm_field_array_int(response_data, UVM_ALL_ON)
            `uvm_field_int(response_received, UVM_ALL_ON)
            `uvm_field_enum(uart_monitor_parse_error_e, parse_error_kind, UVM_ALL_ON)
            `uvm_field_int(monitor_recovered, UVM_ALL_ON)
        `uvm_object_utils_end
        
        function new(string name = "uart_frame_transaction");
            super.new(name);
            data = new[1];
            response_data = new[1];
            parse_error_kind = PARSE_ERROR_NONE;
            monitor_recovered = 0;
        endfunction
        
        // Build command byte
        function void build_cmd();
            cmd = {is_write ? 1'b0 : 1'b1, auto_increment, size, length};
        endfunction
        
        // Calculate and set CRC
        function void calculate_crc();
            logic [7:0] frame_bytes[];
            int byte_count;
            
            // DSIM workaround: Fixed allocation for known single-byte write operations
            // Assume data array always contains exactly 1 element (basic test scenario)
            if (is_write) begin
                byte_count = 6;  // CMD + ADDR(4) + DATA(1)
                frame_bytes = new[6];
                frame_bytes[0] = cmd;
                frame_bytes[1] = addr[7:0];
                frame_bytes[2] = addr[15:8];
                frame_bytes[3] = addr[23:16];
                frame_bytes[4] = addr[31:24];
                frame_bytes[5] = data[0];  // Fixed index (no .size() dependency)
            end else begin
                byte_count = 5;  // CMD + ADDR only for reads
                frame_bytes = new[5];
                frame_bytes[0] = cmd;
                frame_bytes[1] = addr[7:0];
                frame_bytes[2] = addr[15:8];
                frame_bytes[3] = addr[23:16];
                frame_bytes[4] = addr[31:24];
            end
            
            crc = calculate_crc8(frame_bytes, byte_count);
        endfunction
        
        function void post_randomize();
            build_cmd();
            calculate_crc();
            
            // Synchronize frame_data with data array
            // DSIM limitation workaround: Avoid .size() comparisons (LHS/RHS=0 error)
            // Always allocate frame_data and check index bounds instead
            frame_data = new[1];  // Default minimum allocation
            frame_data[0] = 8'h00;
            frame_length = 0;
            
            // Initialize coverage support fields
            target_addr = addr;
            crc_result = crc;
            frame_type = cmd[7:5]; // Extract frame type from command
            
            // Error flags initialized to no error
            parity_error = 1'b0;
            framing_error = 1'b0; 
            timeout_error = 1'b0;
            
            // FIFO levels initialized to empty
            rx_fifo_level = 7'h00;
            tx_fifo_level = 7'h00;
            
            // FSM states initialized  
            parser_state = 3'h0;
            axi_state = 3'h0;
        endfunction
        
    endclass
    
    // AXI transaction item for monitoring
    class axi4_lite_transaction extends uvm_sequence_item;
        logic [31:0] addr;
        logic [31:0] wdata;
        logic [3:0]  wstrb;
        logic [31:0] rdata;
        logic [1:0]  bresp;
        logic [1:0]  rresp;
        bit is_write;
        axi_trans_type_t trans_type;
        axi_trans_type_t trans_kind;  // AXI_WRITE or AXI_READ transaction kind
        
        // Additional fields needed by sequences and coverage
        logic [1:0]  size;           // AXI size field: 00=8bit, 01=16bit, 10=32bit
        bit          expect_error;   // For error injection testing
        
        // Additional fields needed by agents
        realtime timestamp;
        bit completed;
        
        // Aliases for driver/monitor compatibility
        logic [31:0] data;
        logic [1:0] resp;
        logic [3:0] strb;
        
        function void post_randomize();
            // Sync aliased fields
            if (is_write) begin
                data = wdata;
                strb = wstrb;
                resp = bresp;
            end else begin
                data = rdata;
                resp = rresp;
                strb = 4'hF; // Default for read
            end
        endfunction
        
        `uvm_object_utils_begin(axi4_lite_transaction)
            `uvm_field_int(addr, UVM_ALL_ON)
            `uvm_field_int(wdata, UVM_ALL_ON)
            `uvm_field_int(wstrb, UVM_ALL_ON)
            `uvm_field_int(rdata, UVM_ALL_ON)
            `uvm_field_int(bresp, UVM_ALL_ON)
            `uvm_field_int(rresp, UVM_ALL_ON)
            `uvm_field_int(is_write, UVM_ALL_ON)
            `uvm_field_enum(axi_trans_type_t, trans_type, UVM_ALL_ON)
            `uvm_field_real(timestamp, UVM_ALL_ON)
            `uvm_field_int(completed, UVM_ALL_ON)
        `uvm_object_utils_end
        
        function new(string name = "axi4_lite_transaction");
            super.new(name);
        endfunction
    endclass

    // DUT Internal State Transaction for enhanced monitoring
    class dut_internal_transaction extends uvm_sequence_item;
        dut_transaction_type_t transaction_type;
        logic [31:0] data_value;
        logic [31:0] address;
        axi_response_t response;
        string state_info;
        logic [7:0] internal_state;  // Encoded DUT internal state (matches scoreboard expectations)
        logic [7:0] fifo_level;      // FIFO level info
        realtime timestamp;
        
        `uvm_object_utils_begin(dut_internal_transaction)
            `uvm_field_enum(dut_transaction_type_t, transaction_type, UVM_ALL_ON)
            `uvm_field_int(data_value, UVM_ALL_ON)
            `uvm_field_int(address, UVM_ALL_ON) 
            `uvm_field_enum(axi_response_t, response, UVM_ALL_ON)
            `uvm_field_string(state_info, UVM_ALL_ON)
            `uvm_field_int(internal_state, UVM_ALL_ON)
            `uvm_field_int(fifo_level, UVM_ALL_ON)
            `uvm_field_real(timestamp, UVM_ALL_ON)
        `uvm_object_utils_end
        
        function new(string name = "dut_internal_transaction");
            super.new(name);
            timestamp = $realtime;
        endfunction
    endclass
    

    
    // UART AXI4 DUT Transaction Class (QA-2.1 DUT Monitor) 
    class uart_axi4_dut_transaction extends uvm_sequence_item;
        `uvm_object_utils(uart_axi4_dut_transaction)
        
        // Transaction fields
        dut_transaction_type_t transaction_type;
        logic [31:0] address;
        logic [31:0] data_value;
        axi_response_t response;
        string state_info;
        time timestamp;
        
        function new(string name = "uart_axi4_dut_transaction");
            super.new(name);
            timestamp = $time;
        endfunction
    endclass
    
    // Remove the alias since we have actual class definitions now
    // typedef dut_internal_transaction uart_axi4_dut_transaction;
    
    // Alias for configuration class (naming compatibility)
    typedef uart_axi4_env_config uart_axi4_config;

    // Include UVM component files in dependency order  
    // Components are now compiled within the package context
    
    // First include coverage and scoreboard (needed by monitor)
    `include "env/uart_axi4_coverage.sv"
    `include "scoreboard/correlation_engine.sv"     // Phase 3: Correlation Engine integration
    `include "env/uart_axi4_scoreboard.sv"          // Phase 3: Scoreboard with Correlation Engine
    `include "agents/axi4_lite/axi4_lite_monitor.sv"
    `include "components/bridge_status_monitor.sv"
    
    // Then include driver and monitor classes
    `include "agents/uart/uart_driver.sv"
    `include "agents/uart/uart_monitor.sv"
    
    // Then agent definitions
    `include "agents/uart_agent.sv"

    // Loopback support components
    `include "components/uart_uvm_loopback_model.sv"
    
    // Finally environment (when agents are ready)
    `include "env/uart_axi4_env.sv"
    
    // ========================================================================
    // Sequence libraries (need transaction classes to be defined first)
    // ========================================================================
    `include "sequences/uart_reset_seq.sv"     // UVM-compliant DUT reset sequence
    `include "sequences/uart_reset_sequence.sv" // Driver-controlled reset sequence
    `include "sequences/debug_sequences.sv"    // Debug write sequences
    `include "sequences/basic_func_sequence.sv"
    
    // ========================================================================
    // Test files - Production tests only
    // ========================================================================
    `include "tests/uart_axi4_base_test.sv"
    `include "tests/enhanced_uart_axi4_base_test.sv"
    `include "tests/uart_axi4_basic_test.sv"

endpackage