`timescale 1ns / 1ps

//------------------------------------------------------------------------------
// uart_configure_baud_sequence
//------------------------------------------------------------------------------
// Issues a configuration write to program the UART baud divisor via the
// AXIUART register block. This keeps the DUT timing aligned with the UVM
// driver when tests override the baud rate at runtime.
//------------------------------------------------------------------------------
class uart_configure_baud_sequence extends uvm_sequence#(uart_frame_transaction);

    `uvm_object_utils(uart_configure_baud_sequence)

    // Target divisor to program into Register_Block.CONFIG[15:0].
    int unsigned divisor_value;

    // Timeout field value for CONFIG[23:16]. Default keeps the reset value.
    logic [7:0] timeout_field_value = 8'h00;

    // Register address constants (matches Register_Block.sv map).
    localparam logic [31:0] REG_BASE_ADDR = 32'h0000_1000;
    localparam logic [31:0] REG_CONFIG    = REG_BASE_ADDR + 32'h008;

    function new(string name = "uart_configure_baud_sequence");
        super.new(name);
        divisor_value = 0;
    endfunction

    // Utility to clamp the divisor into the supported 1..0xFFFF range.
    protected function logic [15:0] sanitize_divisor(int unsigned value);
        int unsigned candidate;
        logic [15:0] result;

        candidate = (value == 0) ? 1 : value;
        if (candidate > 16'hFFFF) begin
            candidate = 16'hFFFF;
        end

        result = candidate[15:0];
        return result;
    endfunction

    virtual task body();
        uart_frame_transaction req;
        logic [15:0] sanitized_divisor;

        sanitized_divisor = sanitize_divisor(divisor_value);

        `uvm_info(get_type_name(),
            $sformatf("CONFIG divisor request=%0d (0x%0h) sanitized=0x%0h", divisor_value,
                divisor_value[15:0], sanitized_divisor),
            UVM_MEDIUM)

        if ((divisor_value[15:0] !== sanitized_divisor) &&
            (divisor_value > 0) && (divisor_value <= 16'hFFFF)) begin
            `uvm_warning(get_type_name(),
                $sformatf("CONFIG divisor mismatch: requested=0x%0h sanitized=0x%0h",
                    divisor_value[15:0], sanitized_divisor))
        end

        if ((divisor_value <= 0) || (divisor_value > 16'hFFFF)) begin
            `uvm_error(get_type_name(),
                $sformatf("Invalid divisor_value=%0d detected; sanitized to 0x%0h",
                    divisor_value, sanitized_divisor))
        end

        `uvm_info(get_type_name(),
            $sformatf("Programming CONFIG register with divisor=%0d (0x%0h)",
                sanitized_divisor, sanitized_divisor),
            UVM_MEDIUM)

    req = uart_frame_transaction::type_id::create("cfg_write_req");
        if (req == null) begin
            `uvm_fatal(get_type_name(), "Failed to allocate uart_frame_transaction")
        end

        start_item(req);
        req.is_write       = 1'b1;
        req.auto_increment = 1'b0;
        req.size           = 2'b10;      // 32-bit AXI beat
        req.length         = 4'h0;       // Single beat
        req.expect_error   = 1'b0;
        req.addr           = REG_CONFIG;
        req.data           = new[4];
        req.data[0]        = sanitized_divisor[7:0];
        req.data[1]        = sanitized_divisor[15:8];
        req.data[2]        = timeout_field_value; // CONFIG timeout field (bits 23:16)
        req.data[3]        = 8'h00;          // Upper bits reserved
        `uvm_info(get_type_name(),
            $sformatf("CONFIG payload bytes=[0]=0x%02h [1]=0x%02h [2]=0x%02h [3]=0x%02h",
                req.data[0], req.data[1], req.data[2], req.data[3]),
            UVM_MEDIUM)
        req.build_cmd();
        req.calculate_crc();
        finish_item(req);

        if (!req.response_received) begin
            `uvm_error(get_type_name(), "CONFIG write completed without monitor response")
        end else if (req.response_status != STATUS_OK) begin
            `uvm_error(get_type_name(),
                $sformatf("CONFIG write returned STATUS=0x%02X", req.response_status))
        end else begin
            `uvm_info(get_type_name(), "CONFIG write acknowledged by DUT", UVM_LOW)
        end
    endtask

endclass
