`timescale 1ns / 1ps

// UART-AXI4 Bridge Assertions Module
// Contains protocol compliance assertions for verification

module uart_axi4_assertions (
    input  logic       clk,
    input  logic       rst_n,
    
    // UART interface signals
    input  logic       uart_rx,
    input  logic       uart_tx,
    
    // AXI4-Lite interface signals
    input  logic [31:0] axi_awaddr,
    input  logic        axi_awvalid,
    input  logic        axi_awready,
    input  logic [31:0] axi_wdata,
    input  logic [3:0]  axi_wstrb,
    input  logic        axi_wvalid,
    input  logic        axi_wready,
    input  logic [1:0]  axi_bresp,
    input  logic        axi_bvalid,
    input  logic        axi_bready,
    input  logic [31:0] axi_araddr,
    input  logic        axi_arvalid,
    input  logic        axi_arready,
    input  logic [31:0] axi_rdata,
    input  logic [1:0]  axi_rresp,
    input  logic        axi_rvalid,
    input  logic        axi_rready,
    
    // Bridge internal status
    input  logic [2:0]  bridge_state,
    input  logic        frame_complete,
    input  logic        crc_valid
);

    // AXI4-Lite Protocol Assertions
    
    // Write transaction assertions
    property axi_write_addr_stable;
        @(posedge clk) disable iff (!rst_n)
        (axi_awvalid && !axi_awready) |=> $stable(axi_awaddr);
    endproperty
    assert_axi_write_addr_stable: assert property (axi_write_addr_stable)
        else $error("AXI write address must remain stable when AWVALID is asserted but AWREADY is not");
    
    property axi_write_data_stable;
        @(posedge clk) disable iff (!rst_n)
        (axi_wvalid && !axi_wready) |=> ($stable(axi_wdata) && $stable(axi_wstrb));
    endproperty
    assert_axi_write_data_stable: assert property (axi_write_data_stable)
        else $error("AXI write data and strobe must remain stable when WVALID is asserted but WREADY is not");
    
    property axi_write_response_valid;
        @(posedge clk) disable iff (!rst_n)
        (axi_awvalid && axi_awready && axi_wvalid && axi_wready) |-> ##[1:10] axi_bvalid;
    endproperty
    assert_axi_write_response_valid: assert property (axi_write_response_valid)
        else $error("AXI write response must be provided within 10 cycles of write transaction");
    
    // Read transaction assertions
    property axi_read_addr_stable;
        @(posedge clk) disable iff (!rst_n)
        (axi_arvalid && !axi_arready) |=> $stable(axi_araddr);
    endproperty
    assert_axi_read_addr_stable: assert property (axi_read_addr_stable)
        else $error("AXI read address must remain stable when ARVALID is asserted but ARREADY is not");
    
    property axi_read_data_valid;
        @(posedge clk) disable iff (!rst_n)
        (axi_arvalid && axi_arready) |-> ##[1:10] axi_rvalid;
    endproperty
    assert_axi_read_data_valid: assert property (axi_read_data_valid)
        else $error("AXI read data must be provided within 10 cycles of read address");
    
    // UART Protocol Assertions
    
    // UART bit timing assertions (assuming 115200 baud at 50MHz)
    localparam int UART_BIT_CYCLES = 434; // 50MHz / 115200 ≈ 434 cycles per bit
    localparam int UART_BIT_TOL = 22;     // 5% tolerance
    
    logic [15:0] uart_tx_bit_counter;
    logic uart_tx_prev;
    logic uart_tx_edge;
    
    always_ff @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            uart_tx_prev <= 1'b1;
            uart_tx_bit_counter <= 0;
        end else begin
            uart_tx_prev <= uart_tx;
            if (uart_tx != uart_tx_prev) begin
                uart_tx_bit_counter <= 0;
            end else begin
                uart_tx_bit_counter <= uart_tx_bit_counter + 1;
            end
        end
    end
    
    assign uart_tx_edge = (uart_tx != uart_tx_prev);
    
    // UART bit timing check (only check during active transmission)
    property uart_bit_timing;
        @(posedge clk) disable iff (!rst_n)
        (uart_tx_edge && uart_tx_prev == 1'b1) |-> 
        ##[UART_BIT_CYCLES-UART_BIT_TOL:UART_BIT_CYCLES+UART_BIT_TOL] uart_tx_edge;
    endproperty
    // Note: This assertion is commented out as it's very strict and may cause false failures
    // assert_uart_bit_timing: assert property (uart_bit_timing)
    //     else $warning("UART bit timing deviation detected");
    
    // Bridge State Machine Assertions
    
    typedef enum logic [2:0] {
        IDLE        = 3'b000,
        PARSING     = 3'b001,
        PROCESSING  = 3'b010,
        AXI_TRANS   = 3'b011,
        BUILDING    = 3'b100,
        SENDING     = 3'b101,
        ERROR       = 3'b110
    } bridge_state_t;
    
    // State transition assertions
    property valid_state_transitions;
        @(posedge clk) disable iff (!rst_n)
        $onehot(bridge_state);
    endproperty
    assert_valid_state_transitions: assert property (valid_state_transitions)
        else $error("Bridge state must be one-hot encoded");
    
    property frame_crc_check;
        @(posedge clk) disable iff (!rst_n)
        (frame_complete && bridge_state == PROCESSING) |-> crc_valid;
    endproperty
    assert_frame_crc_check: assert property (frame_crc_check)
        else $error("Frame with invalid CRC should not proceed to processing");
    
    // Coverage Properties
    
    // Cover different bridge operations
    cover_read_operation: cover property (
        @(posedge clk) disable iff (!rst_n)
        (bridge_state == AXI_TRANS && axi_arvalid && axi_arready)
    );
    
    cover_write_operation: cover property (
        @(posedge clk) disable iff (!rst_n)
        (bridge_state == AXI_TRANS && axi_awvalid && axi_awready)
    );
    
    cover_error_handling: cover property (
        @(posedge clk) disable iff (!rst_n)
        (bridge_state == ERROR)
    );
    
    cover_crc_error: cover property (
        @(posedge clk) disable iff (!rst_n)
        (frame_complete && !crc_valid)
    );
    
    // Performance monitoring
    logic [31:0] transaction_count;
    logic [31:0] error_count;
    
    always_ff @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            transaction_count <= 0;
            error_count <= 0;
        end else begin
            if ((axi_awvalid && axi_awready) || (axi_arvalid && axi_arready)) begin
                transaction_count <= transaction_count + 1;
            end
            if (bridge_state == ERROR) begin
                error_count <= error_count + 1;
            end
        end
    end

endmodule