`timescale 1ns / 1ps

// UART Monitor for UART-AXI4 Bridge UVM Testbench
class uart_monitor extends uvm_monitor;
    
    `uvm_component_utils(uart_monitor)
    
    // Configuration
    uart_axi4_env_config cfg;
    
    // Virtual interface
    virtual uart_if vif;
    
    // Analysis port for sending collected transactions
    uvm_analysis_port #(uart_frame_transaction) item_collected_port;
    // Alias for environment compatibility
    uvm_analysis_port #(uart_frame_transaction) analysis_port;
    
    // Coverage collection
    uart_axi4_coverage coverage;
    
    // Internal variables
    bit monitor_enabled = 1;
    
    function new(string name = "uart_monitor", uvm_component parent = null);
        super.new(name, parent);
        item_collected_port = new("item_collected_port", this);
        analysis_port = item_collected_port;  // Alias
    endfunction
    
    virtual function void build_phase(uvm_phase phase);
        super.build_phase(phase);
        
        // Get configuration
        if (!uvm_config_db#(uart_axi4_env_config)::get(this, "", "cfg", cfg)) begin
            `uvm_fatal("UART_MONITOR", "Failed to get configuration object")
        end
        
        // Get virtual interface
        if (!uvm_config_db#(virtual uart_if)::get(this, "", "vif", vif)) begin
            `uvm_fatal("UART_MONITOR", "Failed to get virtual interface")
        end
        
        // Get coverage collector
        if (!uvm_config_db#(uart_axi4_coverage)::get(this, "", "coverage", coverage)) begin
            `uvm_info("UART_MONITOR", "Coverage collector not found - coverage disabled", UVM_LOW)
        end
    endfunction
    
    virtual task run_phase(uvm_phase phase);
        fork
            collect_rx_transactions();
            collect_tx_transactions();
        join
    endtask
    
    // Monitor RX path (host to device)
    virtual task collect_rx_transactions();
        uart_frame_transaction tr;
        logic [7:0] collected_bytes[];
        logic [7:0] temp_byte;
        int byte_count;
        bit frame_started = 0;
        
        forever begin
            if (!monitor_enabled) begin
                @(posedge vif.clk);
                continue;
            end
            
            // Wait for start of frame
            wait (vif.uart_rx == 1'b0);
            
            `uvm_info("UART_MONITOR", "RX frame start detected", UVM_DEBUG)
            
            tr = uart_frame_transaction::type_id::create("uart_rx_tr");
            collected_bytes = new[100]; // Max frame size
            byte_count = 0;
            
            // Collect frame bytes
            do begin
                collect_uart_rx_byte(temp_byte);
                collected_bytes[byte_count] = temp_byte;
                byte_count++;
                
                // Check for next byte (timeout-based detection)
                fork : frame_collection
                    begin
                        wait (vif.uart_rx == 1'b0); // Next start bit
                        frame_started = 1;
                    end
                    begin
                        repeat (cfg.byte_time_ns * cfg.clk_freq_hz / 1_000_000_000 * 3) @(posedge vif.clk);
                        frame_started = 0; // Frame ended
                    end
                join_any
                disable frame_collection;
                
            end while (frame_started && byte_count < 100);
            
            // Parse collected frame
            if (parse_rx_frame(collected_bytes, byte_count, tr)) begin
                tr.direction = UART_RX;
                tr.timestamp = $realtime;
                
                `uvm_info("UART_MONITOR", $sformatf("RX Frame: CMD=0x%02X, ADDR=0x%08X, bytes=%0d", 
                          tr.cmd, tr.addr, byte_count), UVM_MEDIUM)
                
                // Send to analysis port
                item_collected_port.write(tr);
                
                // Collect coverage
                if (coverage != null) begin
                    coverage.sample_uart_transaction(tr);
                end
            end else begin
                `uvm_warning("UART_MONITOR", $sformatf("Failed to parse RX frame with %0d bytes", byte_count))
            end
        end
    endtask
    
    // Monitor TX path (device to host)  
    virtual task collect_tx_transactions();
        uart_frame_transaction tr;
        logic [7:0] collected_bytes[];
        logic [7:0] temp_byte;
        int byte_count;
        bit frame_started = 0;
        
        forever begin
            if (!monitor_enabled) begin
                @(posedge vif.clk);
                continue;
            end
            
            // Wait for start of frame
            wait (vif.uart_tx == 1'b0);
            
            `uvm_info("UART_MONITOR", "TX frame start detected", UVM_DEBUG)
            
            tr = uart_frame_transaction::type_id::create("uart_tx_tr");
            collected_bytes = new[100]; // Max frame size
            byte_count = 0;
            
            // Collect frame bytes
            do begin
                collect_uart_tx_byte(temp_byte);
                collected_bytes[byte_count] = temp_byte;
                byte_count++;
                
                // Check for next byte (timeout-based detection)
                fork : tx_frame_collection
                    begin
                        wait (vif.uart_tx == 1'b0); // Next start bit
                        frame_started = 1;
                    end
                    begin
                        repeat (cfg.byte_time_ns * cfg.clk_freq_hz / 1_000_000_000 * 3) @(posedge vif.clk);
                        frame_started = 0; // Frame ended
                    end
                join_any
                disable tx_frame_collection;
                
            end while (frame_started && byte_count < 100);
            
            // Parse collected frame
            if (parse_tx_frame(collected_bytes, byte_count, tr)) begin
                tr.direction = UART_TX;
                tr.timestamp = $realtime;
                
                `uvm_info("UART_MONITOR", $sformatf("TX Frame: STATUS=0x%02X, bytes=%0d", 
                          tr.response_status, byte_count), UVM_MEDIUM)
                
                // Send to analysis port
                item_collected_port.write(tr);
                
                // Collect coverage
                if (coverage != null) begin
                    coverage.sample_uart_response(tr);
                end
            end else begin
                `uvm_warning("UART_MONITOR", $sformatf("Failed to parse TX frame with %0d bytes", byte_count))
            end
        end
    endtask
    
    // Collect single byte from RX line
    virtual task collect_uart_rx_byte(output logic [7:0] data);
        int bit_time_cycles = cfg.clk_freq_hz / cfg.baud_rate;
        int sample_time = bit_time_cycles / 2; // Sample at bit center
        
        // Sample start bit
        repeat (sample_time) @(posedge vif.clk);
        if (vif.uart_rx != 1'b0) begin
            `uvm_warning("UART_MONITOR", "RX start bit not low")
        end
        
        // Sample data bits (LSB first)
        for (int i = 0; i < 8; i++) begin
            repeat (bit_time_cycles) @(posedge vif.clk);
            data[i] = vif.uart_rx;
        end
        
        // Sample stop bit
        repeat (bit_time_cycles) @(posedge vif.clk);
        if (vif.uart_rx != 1'b1) begin
            `uvm_warning("UART_MONITOR", "RX stop bit not high")
        end
        
        `uvm_info("UART_MONITOR", $sformatf("RX byte: 0x%02X", data), UVM_DEBUG)
    endtask
    
    // Collect single byte from TX line
    virtual task collect_uart_tx_byte(output logic [7:0] data);
        int bit_time_cycles = cfg.clk_freq_hz / cfg.baud_rate;
        int sample_time = bit_time_cycles / 2; // Sample at bit center
        
        // Sample start bit
        repeat (sample_time) @(posedge vif.clk);
        if (vif.uart_tx != 1'b0) begin
            `uvm_warning("UART_MONITOR", "TX start bit not low")
        end
        
        // Sample data bits (LSB first)
        for (int i = 0; i < 8; i++) begin
            repeat (bit_time_cycles) @(posedge vif.clk);
            data[i] = vif.uart_tx;
        end
        
        // Sample stop bit
        repeat (bit_time_cycles) @(posedge vif.clk);
        if (vif.uart_tx != 1'b1) begin
            `uvm_warning("UART_MONITOR", "TX stop bit not high")
        end
        
        `uvm_info("UART_MONITOR", $sformatf("TX byte: 0x%02X", data), UVM_DEBUG)
    endtask
    
    // Parse RX frame (host to device)
    virtual function bit parse_rx_frame(logic [7:0] bytes[], int count, uart_frame_transaction tr);
        logic [7:0] calculated_crc;
        
        if (count < 7) return 0; // Minimum frame size
        
        // Check SOF
        if (bytes[0] != SOF_HOST_TO_DEVICE) return 0;
        
        // Extract fields
        tr.cmd = bytes[1];
        tr.addr = {bytes[5], bytes[4], bytes[3], bytes[2]}; // Little-endian
        
        // Extract data for write commands
        if (!tr.cmd[7]) begin // Write command
            int data_bytes = count - 7; // SOF + CMD + ADDR(4) + CRC
            if (data_bytes > 0) begin
                tr.data = new[data_bytes];
                for (int i = 0; i < data_bytes; i++) begin
                    tr.data[i] = bytes[6 + i];
                end
            end
        end
        
        tr.crc = bytes[count - 1];
        
        // Verify CRC
        calculated_crc = calculate_frame_crc(bytes, count - 1);
        tr.crc_valid = (tr.crc == calculated_crc);
        
        if (!tr.crc_valid) begin
            `uvm_warning("UART_MONITOR", $sformatf("CRC mismatch: expected=0x%02X, got=0x%02X", 
                         calculated_crc, tr.crc))
        end
        
        return 1;
    endfunction
    
    // Parse TX frame (device to host)
    virtual function bit parse_tx_frame(logic [7:0] bytes[], int count, uart_frame_transaction tr);
        logic [7:0] calculated_crc;
        
        if (count < 4) return 0; // Minimum response size
        
        // Check SOF
        if (bytes[0] != SOF_DEVICE_TO_HOST) return 0;
        
        // Extract status
        tr.response_status = bytes[1];
        tr.response_received = 1;
        
        // Extract echo back fields for verification
        if (count >= 7) begin
            tr.cmd = bytes[2];
            tr.addr = {bytes[6], bytes[5], bytes[4], bytes[3]};
        end
        
        // Extract response data (for reads with OK status)
        if (count > 8 && tr.response_status == STATUS_OK) begin
            int data_bytes = count - 8; // SOF + STATUS + CMD + ADDR(4) + CRC
            tr.response_data = new[data_bytes];
            for (int i = 0; i < data_bytes; i++) begin
                tr.response_data[i] = bytes[7 + i];
            end
        end
        
        tr.crc = bytes[count - 1];
        
        // Verify CRC
        calculated_crc = calculate_frame_crc(bytes, count - 1);
        tr.crc_valid = (tr.crc == calculated_crc);
        
        return 1;
    endfunction
    
    // Calculate CRC8 for frame verification
    virtual function logic [7:0] calculate_frame_crc(logic [7:0] bytes[], int count);
        logic [7:0] crc = 8'h00;
        
        for (int i = 0; i < count; i++) begin
            crc = crc ^ bytes[i];
            for (int j = 0; j < 8; j++) begin
                if (crc[7]) begin
                    crc = (crc << 1) ^ 8'h07; // CRC8 polynomial
                end else begin
                    crc = crc << 1;
                end
            end
        end
        
        return crc;
    endfunction
    
    // Control functions
    virtual function void enable_monitor();
        monitor_enabled = 1;
        `uvm_info("UART_MONITOR", "Monitor enabled", UVM_LOW)
    endfunction
    
    virtual function void disable_monitor();
        monitor_enabled = 0;
        `uvm_info("UART_MONITOR", "Monitor disabled", UVM_LOW)
    endfunction

endclass